PK   T��Z����6  �R    cirkitFile.json�[s�Ƒ�
��rN����y���YGxm���>h�j��Þm�H�*�ݷ
MٍFw���1�C�B�DVVe]�~Yl���e��t����j}�xC�z�ڴ?U����Vw��z�æ��n���{��Ǉ.�7]���p�2�6��6�2�:��j3�=i�k�W�R-���w�__.��Ԓ����+��������Ұ��Ҳ��ұܞ95���w��vY��ھ�3o�Y�WYi�<k|�j�겵��Ӗ<�߳�-�?g�s%�e�f(X:�L�l���o���o���ף�߀Xo�kU����?u�lS�n�,?�o��j��p�=���p�o��"Tt�L��'��u?p��o1��d�E��4�\���|�E
~�(��[D�[���C67LaG)�0E��A�߁�"8\���A��6I��� �ߞ�E
~{�(��	[D��'l��ߞ�E���'l������{��/���,7��l�uV��\a����)�|���K�2T��Z���ަϊB5�q��������^�⸭hP��(�1^�J�5{�{k�� �����[;��@�o��"��b���-"P�[(��@�o��"���[(��@��x�"?fa�|��( �+|�i���-"P�}'[D���N��@���l���;�"���}'[D���N��@��*Otw[Ք�l}Vԡ�l�Vgu�(����jLAS1F�ɻ��2ۚ2�Mm�sï���h�������ݽ3�q^��tn���-��Pl����B9~�(�-[D��Pl���B�E���Pl���B�E
~�~$b�������<q��#,�
��#��t��SK�՝��JGX:�4X���t���Vw�;(a�B�;�����t�����cu�#,�Z�X��t�g��:���i3�y��5!��UUt���ႎ�z���_�����k�P:�ҩe��]�����tq5�_J�|�˷��C&�����f.�ӬFb�~pp��+����o�|��_b��(�`U��3a_���S]�(��a���|q+X�P	�G`����?hTA`>���'`���,�����������|q�xd�`��7+���~�|����CO͠�f���/����>���}=:�zLu����x��>�����/n[?8����/n���`������~�|招%��G?X>��m�`���,���U��p��#0_�Z�8����/���`��7ڂ��^��^�_x�ƀ�,����f�������|q[6X���G`����?p���#0_�
�8����/n��`���`�g�����|1qX���G`����?p���#0_LV1=�?s+3w�߂C����AT��Z��[��\],8t�������4ľy5���Q�G=X>��T0`���,��b���Q���|1�X��G`��8�?�z�|�)���G=X>��dM`���,��b�&�������|1uX���G`��t
�?tj tn p�����X>��D_`���,��b�2�������|1�X���G`���?�?�|�	����X>��T|`���,��{68�T�c�վ�1��6Yi{���o��m���g�μ�0����3 μ�0�����μ�0����3�μ�0����s�μ�0��\����FG:ν�iy����ϴ��q�s�gZ�舿��3�ot�����~�i�����ϴ��!gs�g���`���3�ot��܆�i�Ө���mx��7:i��'�/-�=/�۟S�}>�������,\Y�LweV>����ʾoU�j[wtp�����0P��N.�a�8�5�5x�Ӊ��n<��^<��N<��p�'�3O�e�F��K�'��}�a>�d=�2��YO���zr�Ϋ�1v<��ă8�N�I�B�6� S�wO<�S��G��$�N$��K<TJ��OWz�Z9�r_dֹ<��4��e�l�v�\��:1��t�t��t�t��t�t��t�t��t�t����\q:�Ӟ&)�:�w��������Z��@Fj�б�ux�r�^6���f��NzX�F�<?�m~�4���7�*�oxD�#����i��@���!	<�$hp��A��u��y� ��lyD9�$H��CT�t�����Jу��#g965�/`�v�\_���#�`L��FM�3�����`��`�%iH�$QQ~��e2��7��7J��G@L Ij�p1�|8��8J�&�AL Ij�lu,a�o�����u�5&�P�D;��`��&�AL�r�aA �	��5̏�$�a��	��5̏�$�a��	��̏�$3Q)�s&�E�	���p]�j�A�	7���GIR��̏�GI���`L0?n`~%)f �1�����q���)����GI��`L�1qܠ8̏[�GI�yu`L0?na~%)��1�����q����6�����Q���#AR�)U0�������v��������Q�b.̏;�GI�{�aL0?�`~%)�M�1�����q����������4����z��a�3B*����Zn��K�U��DX��p+>\*P��$ª��)��R�z�`%�w���0�F�$��A"z=L,�р+���>��^�a4 �J"�{+�z=LDvl}�|H��V�S����U��DX��0e\*P��$���2�-��Ƶ�2�����.������x�O,R�2��m\k.c�2ї-���5�2�G5���-��(A&#�(L��dh���Db"�$C�b��V"�!Z���{Jdt+��Вm�#�[��L��dh�����L��dh�^%���e"�$C�\��VhFLhJL&.�2q�G:��A����B�0�t�	Zff�-Z,R�2q����DhI�6�I�ѭL\&BK2�qo��ne�2Z���{Det+��Вm��*�[��L��dh�]��I2q�-��ƽ�2����DhI�6ѭL\&BK2�q/��n�V+
-W��ˌ�|����DhI�6�͗ѭL\&BK2�1ǀ�ne�2Z����dt+��Вm�� �[��L��dhc�
���e"�$Csp�����e"�$Cs���V&.�%ژEF�2q�-�Ў����X���-Z,R�BɄv�	m%��ˬL\vx�h�W����B� �Y��L��dhc�#���e"�$Cs8��V&.�%ژ�JF�2q�-��ƜZ"�u2q�-����`2����DhI�6�8�ѭL\&BK2�1W��ne�2Z���9�dt+��Вm̝'�[�,Bi>d�2'�9��L��dhc.C���e"�$Cs2��V&.�%ژ[RF�2q�-����"��2q�-���\�2����DhI�6�,�ѭL\&BKi��ΦV���(����Pwm���63m�]�_M��<S�DnڙR&��Δ2��{�����3�L�ʞ)e"��L)��gJ�� =S�D��V2^��N�:W�~��V�+c�S�����cB��X��a�sŀ|0Ɗ�λ�+c�SgA������X�Թ�s[]�O�8W�+���c��9oŶ����̛�eV�U��Y�KUkW���z|�SfJ���,��R�����72�״̔2q��L)�7�Y9S��ьN�)弟I�r�ͤH9�e��I3X���r�Ү���){��/S�e�c*�.[����}aZSs��Mn+s\��PM:km[g�l��(T����*;�{��NT�$)t�RA���]��)^geљ��(K*���ϳ$I9˒{�k�̶��lS۠��.)7����,��o�:���)U������.���eԖ�Q�)�<K���,�r^�Ȭsyf�i��2s�n;C.W^��H�r��$�l$I��.H���=�$)g; E��E���uM��λ,:���}U]�M��7*��?�:���mY��0��:ʬ.|VUm��}ߪ�ն�l�T$I
={�_1��zy������/Ob����Mu��o�QM A;�C�@�v�B���"��]����|	�$H�nH�:�"� 5"� 5"� �R0.�qn�	�Q��.�0�|7��7J��E�&��&�GIR�̇̉�$��\
�	��5̏�$��,�	���u�a~\��8J��Mfa�`~\��8J��M�a�`~\��8J��M b�`~\��8J��MMb�q�70?���v��&�H
n(��̏�$���0�	��̏�$�d_0&�70?���K��`~���8JRLfc��q��(I1y�	7&���q��(I1�	�	��-̏�$Ť0&��0?���8��~`~���8JRL c��q��(Iq�:�	7���ބ�q��(Iq31�	��̏�$�ͫ0&��0?��7K`~�������Gk�Rw�RI��DX�r��-�W	VaU�цZ�T�^%XI�U-GI��R�z�`%�w��u���	Va� ��rA4 �J"���"��Q^#�$XI�U-GI��R�z�`%V�%4BK�U��DX�r��-�W	Va�k�e��K��dh��f�
E]Ba�L�E2��D^"�$Cך��V&��%ڸf^F�2�-��Ƶ�2����DhI�6�a�ѭL$&BK2�q/��ne�1Z���{Jdt+��Вm�#�[��L��dh�����L��dh�^%���e"�$C�\��VhFLhJL&.�2q����DhI�6ѭL\&BK2�q/��ne�2Z���{et+��Вm�[)�[��L��dh�Q���e"�$C����V&.�%ڸgWfa�L\&BK2�qﱌne�2Z���{�et+��Вm�.�[�ՊB�e�2#���L��dh��|���e"�$Cs��V&.�%ژ+AF�2q�-��Ɯ2����DhI�6殐ѭL\&BK2�1��n�L\&BK2�1���ne�2Z���9Qdt+��Вm��"�[��L��dhc��
�$�J&�Y�����e"�$Cs��V&.�%ژ�HF�2q�-���N2����DhI�6梒ѭL\&BK2�1���n�L\&BK2�17��ne�2Z���9�dt+��Вm��&�[��L��dhc�9���e"�$Cs���V(ˇP������eN&.�%ژ�PF�2q�-��Ɯ�2����DhI�6斔ѭL\&BK2�1G��n�L\&BK2�1ק�ne�2Z���9Ket+���R��QѥR�������ǜk�����i������j��R&r�Δ2�Mv���<�3�Ldޞ)e"W�L)٭gJ��G=S�D�R&r>ϵ:��b�w��׹b0�;u��\1�:�t��O:WƊ��+�1V<uJ�\1+�:r��O��8WƊ��5���b�x����b@]	�O�7W�y+���}�g�4.�����<�_�Z��lm���K�r�;�H9��R���J)R��)�ot�ѤH9�gR��w3)R�{�$�/�zz|Ib0����K����=>򕡚t�ڶ�l��YQ�&3NUUUvV����J�r�sE_j_wYnl�x��Eg2W��,�l�*?ϒ$�,K�ɻ��2ۚ2�Mm�zï���h���'�$I9�Ҫ�Te볢nb�Z��s�Q[�F���HBH�r��VΫ��u.�,5M�Rf��mg��ʫ�,IR0,g�C����!I�Yߐ$�k(��.��g�k��v�e�iM�澪��W�K�FIR���,\Y�LweV>����ʾoU�j[w	��$�9˯��?�.���z�\�?/�Pq��i���n��k����z�v�ś��8j����׌G[֘�ц5��z�f��M<:�����Y/�jv9�X1�'���a�xrb�Ή8��Y �;sl��K&hbw��d�����h��$��M�ub�L��q��ɉG�|����%��BNWP�;�u9��i3,l��Vu�͚�
�n����צ�ѽ�]�!���Ͻ?&���NX���p��ϳ�����Ǘ�����<�S ��)���_��űL����0|�]N���<<}�'$�qΠ���O���{�MO%Y^b�"�'�Y:8�G�Aa:����>�(E�V�w�.@�qZ��o���7`z˗����S�����媇�<qqN�ȴ����KAI����%��A^�8T��HB�6�`6�$��\�jF�-MY�N�Js�-Mz<�)?і&=�ٔ�hLS?ٔs��w煙�?9�=�f~��Jn�$L�$N~�����O�Ϊ��_2�W�)��wO(�z_:�`�0;36��1;�'6/j5X~_+6���L 89��"_�_@��6ϴ��0����r���]�����t���z�w��K��78L��GS���I��	���_":f�r�)OgGIfrB2i����/YF���g���E���'.t����^hd`��,)��� �==q4������c>}j�eb#��?w �`v2���g�`v2������<�f�f���7�m����vYݵ�6�}8?�N����y�c �1 s��I���EP�_�� sO_̭e'^b�_̍f|0���5��v���>�p7��� u/��
R7� ����߽L��9> s�ܙ�P~���$.��k���s��H��~��)��n��{Urx���!:�"]B6 �Gv �Os�70Κ6� �ڙ�֐"T� �|���@��`j�(q�@�3�����Hf�o�����Ϟ:���/��ڍ�!= n4���!b /�#vŢ�
.���/�h�,z�ࢭ� W%�iC�N�й,�xX���F^`X�������/���u|���P�Û��(|��\���$)|"t��GB�L��2�p�:Xv����������0`A���~	 �'���������5^�}��D�����/�����lf���˰����)��q����矈���~~��_j<l������.����P��ψ��]�tO.���Fpxw���)�ϒ-Rt�좤��ӌ'��s���(���(RjBI�Q��]���H��;e������l��9y�ROB�-��'5�R�(1�`�����S� RS@	t>�UB �!	�X�����lO�O��'��'�h�C��X
c'�	>�0�����	%G�/�%��/��$��/�e_�8�?��W6Bzt�M&�:�C�'ԁ���*���]Ȩ�~��P���7*�:�&=^�o�r&��._�g��S�'����\`�Ч]�|̡��\��@}�9�@#�Q4����Z���~$
�
}2�*Nʙ�H�C �I�C �K�C NM�C�O���P�I�|�U ��U ��� �1+���{�?�g�;��'��#Y�R��y&�(D��4�	5��$�/^�(D�%vD+�u����k�'��	�q>�k��="�*ƟC-�a��0Dɮ���8vE���ob�_�禬󅃡ױkN����:��!�9Y �qY�bn���[/�ն[������wXn�ˏ�v��N����%��-"��oj����X"���u�lM�E��l
����M�b>��	�<(χ�c�����"Tpml�b�͜�(�P��{1����X9� Xc��k��6#g��\5|5_ư�g�n��	��2T��9�2�I�e�������8 ��/Cŕ4������Wt���#����+l Xf��l�4�笏�sfî��/#p |1_FLY� �b��|1�����esͣ*Ȋi'��uď�"Gډ�b!- ap�|��m�2���e���� o˗8 ޖ/C--���e@ϗ/#p ��|q,�1
��S�|q�?��O-���e�?�� ʗ���O�2���ek�FC���|ډ�b��~�$�x[�|�1���m�2���e�� o� ޖ/C-=���e�������X���Rj�R^�|ŔG`>�%��G`�a�̧��?����|ji��3`�a�����,XX>��X�?,��B? �?����|{�%@���L���Ƹ��/��,���#0�Z�`��`�a���Z����LHh¸.�CxP�J�a�a���+Zy�1*E*`�q"I�@���
�p?�F��x���Y�	LG��@G0��I����a��q�6Z��0LHh¸��Cll@hBB���h��0!�	�B��1��Єq�zTŀ		M7X�u��b���&��A�:�O���W�a�F�-��fOoj�@�(f���((8��'c��(L���ŀ		M�;�u��b���&�[��:DG1`BB�mfh��0!�	�9��Q��Єq{zm	:��p|J$T F��(L�Q�u��b���&�?�C�B1�J1t�bГ/��		M7ۢu��S���&���:D�)`BB�M�h��0!�	�m��q
��Єqs9Z��8LHh¸1�C��S���&����:D�)`BBƄh��0!�	�ǉ���2�o��e�Q)|�|�|�:l���𐺑���#40�j �Xt&$4aL-��!:��0�EA�ŀ		MS��u��b���&��h�:t�(LHhJ�Ct&$4aL��!:��0�,B���		M,�u�[���&�ɡ�:�oχ��G�)�8t�&$4aLʅ�!:N�0&C���		M���u��S���&����:��8LHh��Ct�&$4aL���!:N�9�gGc*U�x�y��x��6Yi{���o��m���9��Qę���μ��u����3�%M�y�(����GIJg�?J.:��QRй��6@�����+�k����
�Z������v8>�l� �%���+����8>`k� �%���+�k��#��
�Z��P��m�����n���8>�g��S��rh���Z�!����!�H�~�gά=�)n|�������'B��5S��,����f�;�pR�?�oR�?�n�,�IpĶs��#��8�X���;b�{�s'�ϕ76p=�k�W�j�Yk�:�e�gE���8UUU�Y��#�p��$�;rN߄���/���,7���ʢ3�+LQ�T6E�ϠK�N�{�k�̶��lS��-¯���h�����r�I�Դ�F�UM���gE��F24�u�(���
WMA3�ĥ���y��"��噥�����ٺ��\yujl"������Ot���?�J��D(��=�����|溦�l�]V�ք뫪�z�;u�fMXG��#5k��mY��0��:ʬ.|VUm��}ߪ�ն���D(I�:���z�$f�.��e��x��"��x��"j,V����]����걑��%�����e�*ݯᅆ�oh��Fuhi��a��z��������������0�3��;L�#t��	������>�b<=3ܐ���nH�{7����R*�ކw:_}���`�{74ymu�)+�
j�m�}Ӕ�6�w�bI�z��P*���PD�<<���t�1��}m{e�v����1�C]�"Kєegv%뮩��YgT�f}>{0,�QN������{k��fd�9*�̾�:����Ē�b~��ǻn��rw��%\��8�d�90�L���c8ڃ��wK�a��1��Z&�=�C�"��X��)�Ƅ9�����Zc����8Cbd����cE�\EL�LbL�]�D�#E�b*�qF�x�'l+���Ĉ^b��I儔cE艆4qh���w���������Y�DMJ��>�r���<�f��a6�\�c�8m�gv�#��˦�ǲ��#@9���蘻.XD�G� �, �rc =��r���ų r���]�Vuwc�����m�b3vp�?\��K�p�Ɨ��%=��.����R>�T<\*ƗʇK��=��_�>я������L�p͌���kv��x�ȥG�G$>j����OC�oC����.�Q�4V&=*���ԏ��èau{�|f���~��]�o��kU��&�Z_�NWmˬ=���n{]�Z�1�^�u�[+�y���!�y��LuE�-ʬ�M�iSZݘ�U!����ެξn��U]k������kڬp��j�ݻ�Е�X"oo\�)ݍ-��	�o�~��w��=��)�xN�pw��S�'/r��j[���v���m��n�}��.���#|���fu�Cx���}�=^�^�X�~����ϿW�p>ޭ�"�����O��&�]����.\��6[ݯ�����6�\m�v�fP�U���>�U����6� �{F�?���@PB�u�]���#Oōu�C��U��«�O��F��	�������
_k�}���rcL�����K����O�����~[�5;AI��׋�f�T;�E��)~�f�in��o��V߸�¨�?����6�j�E��K}��t�vU�:7���<8Q��X�}m�.
7Q �Q�rNM��	OWN�$���:����롊���}��sun�>�H���{���u���\�я�B���jC1eoBT����^���8�E�����e,P�S$�܆7u/y[�'W���H��w$9=��D1��f��L��� 9q}�Z�b�V����/ۏ�j��LtcnL��G\�A�	_���<wי��mpHv��Ҹ.h�nʬ1.�H:8}=D�emMgt���J�*M҄IZ��.���&���?v0��Ec�=�� jO|P�C-�H�+��"�K�=J�E/��z��]���j͍ۿ��^p�������_��]���S�P^�Lڡ�ǁ�
�S��9��b�ow
R_�e�>��օ�ɝyBp�U,%���T��U,N\�Y���;U�u���%M�n����v�=㢂��W��Qy��[�d9}B�J��C[�T.O����,n��C�=���C#�sm�=gR�V��wY�l躄BYUu��n�NW��Kt&	Ӷ������1�ҩ�(�����(o�5�?�%��ae^VaI�։
Ӕ?)�J�),���C�=����Dg���S?��u__�a������jۅwy{���o��m�C��*���������fn{s��W�z��n�c?��u��|��'�gy����'Å�]/��Շo�䷫�V�w�~z�pS�����?l���oַ�����a�'���9��O���C�����<���:)>�L�?]}F�������n����tG�~���h�J����ͪ�=�_�� ��&ϋ�/(� �9S�μ1!Ry^��1��uV�V2k)���u�S_U6�
���60i����Ë������z��\����]���?��ew�������g[�������p��_>t]��J�Z����j�uџ]5��\������R���������Mh3�&�Q�-oB�\����M^�	$-{EN���mw�W�f���]��Տ���AS<��\�����b�P�.��c�کX��x�Ɔx�4./D�uҺ�WT��ڴWw�?V�_6�W_��}�CetquX���g����/���s����[��©�&��F�����*X}NZ�������v������cl��ɔ���_�p�:�/��Ku~Ѹۨ����yh��UtM:��F�<��ܹ\�6�����s�ڿڍ/�T��k� HF������O��}vU��Ϻ�٬+m�y��̕�
_���,�>{����V���c�k��S�����Dy6Q�N�Gi�Ty0?:*��nH_���g���YqC1�&M�IS)��2I�ؠvS����t��Ȝ�Y��b#c:^ldKǋ��9^llIǋ��x��/6����Fvt�؁�D�;:^�Ў&Ԧ������z��ݙ�+'����]�QiG����:6C:w�ܰ�����s�_߶�����CC�v������ݶy�vq�v�j���ƺ��mV�gV�.+�i2��ծ({7��~��\��?��o����ke;�gu�]fm�3�>��\�l�7�+��{���guY�e�g�wq�@EYYEV�}h�Ke���~�������;[�VϵMf���Jӹ�qښmw/x���?wQ���}l|���w�����&4wmn�l۠�:��U�ĵ^{e�R5͞*��6���O��gRJS�p[�>�6t�4�YQyZ�.]hT�K������{NӶ����3�kZ���i��.k��"w:x���Cu�v�!Px��v}�������w}7H|����͛��n=��������oכ�Wm������zM�V��~u����Ճ�3yct�M֙����jBg�WM��v��|cK�J�Y��r>�
=��1MS�yg�>fa]�5&�� ��*�k)lVQ_%�J;ia��U���_PӡJtEz�Ee�9ca��׷�׫���~�����/o��]]�ۿ]��]�c�q��rK_��6���v}��xw�ݳ7�t��������������M����]{����v��n�f;��Cਮ;����ۧ��M�@��禈k�ʸ.�ҍsEQ��d�Y��no�R��s���>-|X����?e�R��݊��"��o:�ί���c�<DD�u ��ohX�>�^~��)L9l��i�n�E	.���C�?���0y�j��Q!^�a����c_|LbQ5���OK���t��?���~�����u׿D�Ut0��M��`NA�����
t�n���kO�J�\?��T?����;���zu���ھd�Z�vW����6^����ǿ��.�{�����enճe�����b4Qlo=Lr��53�c��-B��}㠢��k�4:a�d`c�����k<�֋M}��b�ƓV,���q����맬⒴P�8�2q�4�x���u�>�Ag�
~��q��b.]�;��b���d	�ᒼX������	��mE�	�K�&�@M� O��	D�A��1��&0��~��!�;j�>cC3�`M��HC�L��l��(0m梆�+\Ww��������#���٦�"ֹئ���>�U,�}ڮ8Q���AZ�'Q;8+\�ʵ<��%ņ��X9w���3��T]��Sf+�`������D>+G��7EJ�m0��#�C4�4�2��:���/���ݩS-ͨ�볃��z�v����`���TB���g�:� -š�$7 3X�v0�2�vf�X�G!��Ǹ�q�)��]�=U{�\����B��0Ty��B�ڙQ��gi�DE� ���ʵ���!߫٩����r=�q��g0i9dE&�����5��&$wj�`ҊeT7�!A��r]�.��B̩��yzƀ[�&O
U�f�sF4���r=��ArK3��kMH�.)��Ǉ8�ƨ��3��ݢ����`��TR�5Gc�Z��Îɸ���oss�C��R���ϙ�
�m;�;׀���T�ʛǌ��c_~�I-6��{(v0}�[�17�=�|܅˻f�"���l�yJGz�.|���O�?s���=����Di���%�q�A7�8�R�N��bKB��j�l(�Xb��B��ˊ/X v�>.9B�;sv����D?����S�)�a���OV��92��x��DGXU]�p!����iyv��a<1;��9f<��
}Y�D�itє=�x���$�w"gz�=v��S�b/��hbm�~���bOy��L(��/�M-K��9{)��r�w9��2i.��hbIҧ�zN�Tsq}�Zx㔶i*�#A�rv[�e��f�x�`���D���3��L��tق����ًG����\�O2��b�D3�wpEb�Tc�qZ64���m,���V.�1:(V�OǗ�(��Yr[��@c[0��rْȘ�%�Xʃ�/�{${g�$��2��}u{���?�������M������t�Vw�ۯ�����Ǵ�}m��f���f���٬><l�_���PK   T��Z����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   T��Zo�>��q  �q  /   images/2cd737db-51bc-41eb-8762-f3273c40eae5.png =@¿�PNG

   IHDR   d   �   J���   	pHYs  �X  �X{�M   tEXtSoftware ezgif.com�óX   5tEXtComment Converted with ezgif.com SVG to PNG converter,)�#  qIDATx���d�u�+wuu���9�LO�   $ DҴ��l�Ғ�//�����o˖,��%�f	H�� #@�<��9��t��s.�}^������*LWx�{O>��+�/�xF�`�5Ci��� ��ɂpE����0�(M� ~>�ؼ�Ϡ��E�h�slyh�lz�k�.����ޏa~?.�7*f$c躴W���8��F����kX'L�{�������������;��|O�ԏ�G��Iy�7�r��f�l�)��ϔ��_��R��zmU���˶ғgsy��YX�&ē�Af\|�j��,������XC�����B����c����
�k߅��,�๸zb$?wD|roS�r�$��%����׭�u���fHL��e>��0�w����q�W'3�����/��'�A�s&)+c1fL�0�y�����xP1�O�^j���-�^�^�1C�ɰ�q���K�pq�mȘ��r�H�z�Ɉ�3��e�:��U/��_R�|U�J��g?ٿT/a�}��=�^�׻�U��;��ں��>����Q8Jl�%���3����9�}`4
�JSN��蜼a&���~���� �qj5Rg𚚘�"dN���T���yo�x@�K�m��~u�fܱ��F�շ��jZj2��.M}�W̐{|���O�aځ��]?����m���w��+������돖s$f�݊P]����=����A�g䷅�Иn/1���V�O��߁�����͙MbN'(ok]g�V!.��%�7���PO99vje��M娭.��T&��&����1_XM��T&�Z�u7��²����Ȍ<��;]�/�^��_��n���y[gF��~��a��g�`�u,�!$��8��b��� �V3b���J�*��ho��4�W��^Ĥ'R ���4�Z�X�U�V�nW9��¸��]�82�dL��Ɂ2G	l6�.�z�Q��.��'W���D0���w�_B���������m��� oc�$�}B'�{��[�j��>���7�N����oe{�!(ťQ��/m�+a�P8_(
���:~9�O����5ÙV�հ�5msAL��KHnv�Q��t�l�� ��UR��1��.�t�Ӭt��V��`8F{U%&� CA_�41,c�g���/�h��"�X��AӮ���E���A%��"�_S>�&u8���ΐ{�k�z�q���i�����-�f�ɑIܮd�_�qkj]��d����"FYi)�������I��9,-�J�8�N�J&10�E8�+��E�(ä���9�X�xnIf�[�a�K����+aK�`���]�h/c:C��L[ZfDf|S�6/�.�������'S��T��<"Ay�����>̏#�b^¼���7C�PL##����`�8�ל�L)�a��d�d��yJV9�������p����_������H0Z�����[�������Zh4/�x�������TF�\r��p�e��lƺ:7�?�+�I=�'��=WE4����ai)�^�xj��e��D2�٫a��ӞP�?>'
��M,a8��A�#�Jǐ�]��8����A�uU��K����ك!�?�(�[��,8�+��8�N��[���Ħ�e�+�2��,��U�eQ�>y�,�͍5x��E�è0����@�W���U.~|c���*�Q���:�M�R^���"C2�)dm�I`6�5Q8��=~�vZ�J�a��#�?�}.4��3i��
Z� ��hi־>Z�E�9�ECi���9�F�/d�k!Ys1�a(� �l�P�L��T\-5�ƹ(��4*��̱83�3?���4e��$�:sB&�@ځ��2�sFe�L��,N�"ڮ�Z�I�.���nRք��8�a��	dсH%����Vem��]�z��M81<Y�3�$���i~���	���xlp>eyݿ���	*��u@�o-��S�#�P����U����ؤO�0���2Md�PVQU}7��~ e�b��Rq\<�.�~S��ȴs�V��*$��]��OO]Ƒ�qaC�5e�p�,�V�,�A3}�@>.ǂ�妭��ýsT�0S���3^�8�������Ճ7.�''/#O�t�.���!l�p#�l�[Mv-ҞLFP���>��z�S+�S�Ȑ�Qgv��(�6�:@���ذ�$�a\�tX�y��'����E�ꮀ�j��3.���|D�������[�aH����7:E� =�DzQ_��1b�9�ڱ�DF�X�8^�Ua��nU�e�HT_ ��U,c^�����(�����dZ9�a�[6���5X��~d2i���V�l��]"�↨�Dj��S�+�4�n�����_�4��f����m];p��	�	t�&#qE����كjFT�m����;wh��xbY��E��*Q_��\ex�^�>7�ya��S�6�`]W��w8J�?��/�]�82��2a��F	J���e���g�+��p5v�� d�zQ�әt��h�%�ؾ]�ӈP(�hTcHYY�_�hjߊ����zTK3����VR.�������.�(�b2��J��s�$��(�?��4�܍߹k��c��b������D�j��� ���h�C1�4Ӑ��(u�p$�Q�ʫܕ�(��Qj[V�y�Qf�b���Q�j���)T��g��t�θ���lu�ԘS�ȋJ0>�*�/.Y�7��ۡ��P�IV��h�L�+/E��G=�~�6��7�T�dX�7�Ջ,�3�7S�E�dõ05x��� >��M�EgS޹2�hքx&��o�����3�΀w!��t^���"��b|��G�P]ی��!�I�ӱX�hѼ�����_oǀ�����:3�ş������_|�nL�cP4-1��x��t2#J��,�d`��sIu�O���Y����2â�-��T0U�`^Q�~������?��K$k��2m�{��a�N7***�����0����d�R�f[���K��8~��X��.Tմ�>?.����e9��@M��><0����(�a������>�?P�Դ�U����R�5)�8}ދP$�&�҄��sJ6�d�(�:'�;�Y"J�_��:0��s�BPD}\Mʛ��ٿ��s�S��B�������h]w;*�u��o�^�Ao��Nq9�1r��I�<8{��ܝD<�DU\}G?$'�/}�&W9��=7(k"%v�����	���,�a�-�9J]��o�5s��S�B|#Ô�+�n�¿Ӵ�Nxb3��i�N���X<m ��/���_�f�_��d���2�_SVz���jS>�7��x83
�i8�er��X�#��I�Y9���4>@�/��0eՏ�,�h��\�_w�6��K���G�����sd����Y���T�[݁���3*O�xLZ)�ц������w�@\��i왨[����ʴ���B	��(5*�9Yۅ�����e�,t
9	��4�9)98��%��d����-x��i7FR�c���|{0ZQ�O�%��y^�d�Z��YA �U�m��o2%�H8Eg���=��Wˋ���-jA�F&٠��dm�|ҫ��Z+�rt��&��{�*%��)�t�?�s3j��sT�����R\q��.%Jq�P��;�2�GQdY+Sf,�1+�������VL��$�v����o߉py���rL�i�J����������[�8��r��|d�|�����&�n[638RjE|F����~�,���\/���%��>����)�rb!N&�^h����>Ҹa���>�jʚ�E��u�ߜ�~w3t�)6�s��
;��nI�&k�B+�[���s;�x��E�$G��\�tg�E�9�Xd�p�k�7�9�:sR�7c�xƦ���C9Y�<t�L��R��4�(TY�m�d�ErzlJnX����vqE�ߧM�¤��_
�CjcU��?��)�Z��F���9e8��I&����7"�Ί��O�4d���$�6%�ϔ����	�OŲ����+&q�ÏjG�� �Xg�6�$� OZ;�<V�0�̐��Ϣ���6��z�A˖�sX��\������|u�]��_��0'���qiZ��8��'��cq�"�L�T�����PT�}�����1�D-��XY�WN2N�jK���FG��r�:�co�/�k$<��MQ��ϸFqWMk�<��n1{#!�N����~|�ӆ��*rw[=�{�,.M������X��;�� �~�y�zK������oܲ����F����qyҏW����Y&��@����{v������僸��N��85�A��&"1��}�o�/���fū��3.{�V�����\3��V���h���^u��@5�4~��[��v�GQQ�CBJw�{������h�C��]� nq&��/���	���i��۾�D��79�暑)b~d�ZY��~�����=r'��{=~��ױ�wX�m�b8o��R~_�syXf�ya?��7I�W���1���{qcg~���xJ�<�$*����AyΕ�-��/Wҗn؈�/���=nSף�Ģ���ٖ3��W׿��Yy�!���,E�����:�АQ�����f�28��V�d�[8��p�)J��y��$ �ު��CD"��f�Z�vW���Vly
���Z%F1�XC1u��v�W8�~����~���Ͻ�?�м�U�A��P^b������$s	�e���G���W�ƍj�S�Xc�I�RE�l����-Aյ�9vQ�X_
+q�xۋg����Ŕ 6f���5�5�J��+��ɘOo_��)�w�����0Z�|%%�������(--�PJ{�lۋ��!�1$g\�4�*�E1f���uO���Ҳ*T��(3*���+��y�6T)낡���hQ~2O��H�s�"���f5��ֹ%>ƙ��ۋ_�Y+����n���*�'<���5�2591(.�&X�����~�
����qD����FYi7�5���ʛ���j����|�<K���	��*�98Ԕ/U�iH�&�Zy4�L��V�(#*'�[��i&��Ab��E��ň�AQ'��VM����h0*L�\׽f*�?���N1��Мd_��D�~����R>��5�Z-����~"q�,�����*��G�Y��W	�=ј�r��o\]ĕ�����#%�ۧ�j����\������Nq�;�+�k�^;x!��<b� ���w��FD�w���j��!�SJ!�S��&���p�\r��b�0r�8��F���p �̿P�Œ�}]��'�L�;�O�O^: E��2���s*��s��)3����3�"��R���aa�o=��X2�� !#�X陚r;B�c��ӭUZg��/J���~�������ij6]ۂK!~Ef߽�M�	���iF����i=ʕ�ŕ����F�O�r�!<(����F���Sr��Oѽ�>�W��g�TO�����x5� "��`�(k�ܸkj\��{��o�(�$z��#�����"���	qEP��z���^%�cx�L!�c�siǘ�SǑ���Z3��Fÿ�c��C��߾ye����ڎ�^�>�<:�߆R��2��q��k8?>�wc������?c��<���H�qT�[`4[�c�7��kq:^��!j�ݥV{?���I�|�
�y�mE���H��6J���P_%��R�E��ӣ^�I��uI����iҲ)��7u4���J�E��9�X��Z�TsL�����E�N�@V%�I��}�d���^�Ӝ=��(.����Yh?O�=��d	�z�[��'�%�8�<���6Yzz�KKG�2�ej%����Ĳ�P���A�S'���ރ?{�Z}�/n݊�z��]��XU���l�§w����]|lC��q>ea���rO_T&/E�s�{���|nZm\!��1X|'�Do��BAԍ���K9]�ɚfĸf8	���(oG�xnM�C�dM>R|G��4?���Qu#&���o]�v�Pщc ��{{ڕ?��ev�I�$Q��k�'��`��W^;$���߾s��MW��c��i7���tʹ�J-5;�8�k��eD%�0A�8��R p����o��]��z���ӆ���W�ʭĘ[�K'�֮&1>�R��M�P��s�����Y�WOH9�sA7z*�7�7����S����,~A9t�Q"�̸A���UI��Jaڔ����٩^|�|/+����m�老C�4��k���"�K6�:��p�iW��\�N�0���C9��h4gR��aNTR�OVc𬴰H\z���Qlo�뉦0���p���X\|!��_}�Q1|S1�޴	�����ӧ��W�Пb��B���t�)����z��t�*��2٣9��8Y<h�=�[4ZSb���F���/����h`�ɋg�Dw��Dx�| ������и��ƊM2�0]���0=� ������_�}5E''��G��C$�������防×��rv�����CI���58�(�_��w��>�DG�&Եl��dE�;���c2�L4%�󚼤���^F8��)�z� ���&��"����B�]��7���C�B��T��E5{��
e�"U�_�|�I��k�Veб�V��:����]Ės��Do��f��dF�-�O�&�u����=���XQ�Z�6m���'0��⥐V�M��*&�8X�z-g!e1����eI�?�m�]��[׈N�2])}Zd��cJ�3,O���k59�3�&#����5����7���/���^aƎۿ���v�DZ�������a0e�ج{����^�6u�m͍�E�H$��Q�����tm�7���ވ1�@��fl�D,��w��J�+���l��z�2��wN������)�͕I��*�m����������X[�߭�"�=(1FCQԖ;��c���þs�U�C��P�����TJ����醵X۽M��4.'����R�4Xp�vZ��bkV0:epV���nB�)���8hgl^)���Pj���ޡ���,:���[E$/r��Y��>���������Z����YPJ������|��볜��o�$� ��{q��p[������ee9Y%��c�*��
K�%�󘲜��l�PԠ�ݥ%�፼��UWUʿ��*yA1�Wv�Fc�	Ix�p�����7��VL������(���>"����S�L\񅋹�tZ3|�[��Y/��˹�C�tG�vx�.�}������`�
&F.a2�G0kE��{]+�V���a�����lZL��3n�\8�r�ҙ�bJ��Ă��،o+S���ݿN5Y�"a�N:$�&2�7ٰ
���}cH�,�eL:���u"����զ@C�n�	fd�Ǫ�{�N��������^�V�����*�W���ɬ��Š��Mba\�R�3�N�����7 !��:�^R������bV��ad�^J�+�`m�m�P/W>��6x��Mh�ڦĔ�M�Us��>�]T�i�Y�`*����ѳo!���~�t�����C����*1.-ګ�9�yCb����c8�����ء�'���)�c8E�3LQ��h����<?���=�L3;y��V�0�!�vI�O���L\Fe��0蹂��^<�U�����qb"cŭ�Q4�	��i3�\�9��.^�=e9+Mh�9�"�!�U�j�����տ7����\��l�t��X8��0j͞�ՋY�+rU}�.k8e���f)/]4���E��O(��:�� 8;g(WC�_ж���c��C'�F*q(Z�cN�x,7U�=}�	��?`�]�ȟ]��YJ����\�!�+��=��4��X��w���R�%#܎Y%�T���EKQhCX���O��i��.��u�Y�x_ؽAV
����B\����C/��T� 4O���h�Ӝ�N{ m��0�E���.�J�ˌ�	�3��+qE9B�T68�㯝x_��}��-����Eh���G�Lɂ�^�<�BWU%j6�d�"�����i�����n�p�Gz�j��� ��w0��8ӥ�E��sm�m�bE�g�g���I_�KKB1UeNĶ���a�'�W�Њ�Ez��v��+n�U����ӽ�pWJuű�	iN1���1Nhf
!�E� <ӏ�ou,^��� !�i6�5o��H(?�v�B{�^:t5�(�*϶��|[�!y�#b��Sk[i��'�i��б�&ɏPtf3�9�&L���_��I�ŗ0�:c�Ç��jl����؈HD�bd�Yk�n���=�3�r����Şz�rGs��CҴ�8o��������-�MR���֊���d�bc���6�uXR�"���K2��'r��,b����]�ޟ�K%�Y8A��o�;��3�;)3�=���n߈Dx������`$�eh�؂�u7�F�P���T�;D���OC���K��˥�A]�͂��0���Ӳ�J$a�|�� O��f�U �6d
���2��ě������]�]���|�Y�׭�4��C�&�mz��rg�nu�C�c��vIg������qɂ�r���Ȓ�<�9��]�B��`�=��$�&)l��BQϝȸ�VU!�bN%u��*ڱ���^ZC�K�B׮}��pZިt�1�n��5ɰ(�b�7o�,���К?Y*�r�\Y!�&�����7%��X��C�*"�-���C��ݒCg��rǽ��$�2@�bQ6�t�XGt(�}����,��)�3ׯG�R��!TF��RY��i�k�����_gBk@ �Ƽ�@��z�ח�"�P��� �A0�A$G�g�ZC8;�Q�����d� ����a�e0,�(T��7P%f�d�:�d�1rJひy9�2>�OO�j�35I�g�߫VL���@q�ʹ~I�2�lf�~8��׹E���\JWcؖA���6�D���S�b�(	�@]�"j�N[��;�o�,<��1<wb��E��AS�z��:�^\؋S�2��b��h���	�̿|�&��Tc���A,=����<j��H�ܪV_D�����B������!E�>��-x��9��bI�r*\8(J�r��i��+�qbԏP2+zc4�P�c ���}�e2�u�RY�FI��Ա=�R��狪kJW�ҝ��'����cM�w�N'*�|E�׺n�,q:�"v
�ѡ��?��_�T>DDq�D�o�����G��D�	'1|i/����R�Uۘ{��K�����s���B2�ŗ����L��F�P��TΣ?��Иbʬ��Z��U|�y�i1��������q��f\�g� r�R<�Y����JN[�6wwng�Ą��6��O���0)E<*�n��j���ܜGu��S.�JY[g�#MF\
��S)Ԋ���\��J��E���F�m �O���&8�͢�~_ޏ�}V�T��̎���������������P�I����9��:��QD�c-��ڍW/��̌��X�L�V����9��^���������+-xl��D���lbQ�~eĀs>,9(2���wYQ���t��:[���98G��ޅ̒"P:�յ?�aC�#���
��/�)�}<~�$Ք|�=\TFC���PրoxZ���6�_R��"��������U0L��1DS*�*�u�ƜU�/ˬ�� E1e����<���mk��)e���ӂ�λ�51�t;��J�e��Q^�Mq#?��u{O��u�c� U�3rGYu�Dte�u0Y�72��k��g�6�-��$�D<P ���"cJ��`��'˟XֹX��l��
u|�7u��b<`K5��`�&q^&�w�����)	�Lfl˴`[��.�hΈp�
�h���e$��iv�a͔�e�:򕔽��Q��2��t!�b��,e(svA_�LR�$K+��4�b�����QKiC��4��D-���q,w�Vu�f{]����)�({�r��G�asNnOF����=c^|9�|���hɂ�=��dMI�bFYok������~{���옪6^���W8N�l-W>;�|+�K��2exH���C�,�Ȝ�!:��>�L�O�3�ɔN(g�F!+��2HEF\���=W��
�������sq��e-q�7�[�#��ҥV�n�u��h��ԗ9LdK����倧L��1��a����2�D�dRQ�Ux���t��b�m�W��fK�&��1�8��)�E��L��R���3B�E��{�v�b[y��*e�*���rh�c����×�������M�T��hi�(u�Eɮ`m ����OH+v�]��!��Sk:�W+�L�R�{bnN&�G  ��҂�]h/t�f7��U�Õ#�4�嬕���&p�o���+G�1�)~�=���ʱ~���j�fC,��ӯ�y���p19ϦO���B��AX�a�n�)+�
3FKQ/,=��Qq��j!�Eq��:�^T�%�G6��UE���u��s��z,�z�#�q�7[��ժl�ڀu���>>c,�C����P��7�m��h����Ƕ*#���"FUZ�r��vJ)�{���U�Ol��~�X�)��9g�G2���R=��(��zh<�����V�U���uk�N���X|����Z������-[$V��&[����#�+Gwc6����_ ������ �&���x+Z5�-Z�6��в�5��������Z���k�.Jӛ2a$��ݛ���=p�l5���Q��%��KP�&���~�f1�mW���rJG~e��a����yv{#�\-��b�k��g����=un��͛��ы���S����]Ꙕ?���+����]����8�*�*�p��eƬR�.�o4[��=��I�,�b�Ty�~�����ֶ
��3�/�Đ[:�
�ۦ�ei��C�DH�'g�X,���aͦ0�G��Z��5c"
�3�����	\cv���h���h(l�\q�E'��4��R��$:��+%reT��b�7[$�+�My��P]Qt���!_�k�����ա5�O�:�p�[�L�/!��FB@�<3�7I��:5��q<���@L���K)��I1Eo�  ��ҙ����V����Dc�g�W=�U1٬<�d������5�2�l_.����b�I���L֢a`T�q&��9�,$��Br.��d�h�ٞ1���J�psG�o�;�?�����$j:� �S/�hV�'gf�&+�c�,��ݨp*g�l���
I)�=t� �$�ZC��QȦJF7�z�VJ>EY�J�&�N{��u�64��m��14(shp�t�@ ��b���i�6�J'�U�	�T��H<������Ԭ�xl�RXJ�i	��:W?���粪s�&�^���\�S�	ß��n��/U���èm�H/1�9̬W�{H�l�\x C�R��Q�B(9�,:6���)E��B述��.��pK�Q�����XSf��_V�.���L0�+O�f�&�#��Y/ȝ-��$6��)e�D� �a��� Y��[ެ��\,��!���RDLd���x��blԤ������;�+�d;Z���O0�Ƌ�Zt��`>���N���+��{�w�U��*ڷ�,r��W��=�mV�� �.�J�Mf%�|�%���i�(X�u33��B1B4� �/�h�w���d��WYd���Bf��b���#{����DFrKβ�������I"K`�����\ȿ{�0o�6?If�t��z�g�S���JY\�����<�@���ʷr�"E�86�i��~Ά.�������Vt�chS�#��2帐l`��:+�Ӊ��q�I��`x�d�^�թ�,3���o�>aN�Ъ1E�p*�౦�u���hn^�$�q���x�~,���C���G���$HC3+��8w�/SXg���}1���66�*���8L�D�������7��6���5űYD�s�l�Q0����.'����b˼"Kj�a�K/��H��ł�CO�c�ֺ���H���z��ڗ����T���͢T��V���4�
����^�+l��0��"�0�8�79�(wYar�Z���A� W������_�,ZƐf.��c��7�U(�����3��CgD�)�I�z�V�����rnqxQ[����us<V�L�Z�v2M��2«���˩q�qD����$����^��a��t$��LY�W1���a��J�h4��#�)����<�i1�!�>ZE���Q��#=�!�:ϼ��~�J���&��X�IӮ�¡�Щ%�� lo���8�tH9>�c���R�C߆�FҀ�L�pp�_���:��<
gU�����>�9�*����`C1�S��n���g[�|�-�}�e�q�b��o�?5�g��M���[1|r[w��|.�1f'�MY-O䃛S-Ҽ�Ǉu��y�b�G����H��^<X9��5%�q�?AYy�Е��c�]H��\L�q*^>U(Ǳ��GS�:�7�G8,F%YL�ߎw`�ĳx9\�Hƨ����۔�4]��KoD$kn>Ih����[�(�0K	e�_���]j-u:މ�/;���ŭ�V��H�=��b��$Ƶ.��a�=��5�	3_H�n���ـ���1yH�QR�2�P�- ���L�(����i�W��i3�A�P"��@���!�o^\���<�Z]����%���XY��"�2����R[�%�+`�N����1I�V�)��!�҈7ϭ�~p�@1UX�rg�������)�e�]���d�3�5(��8���L�_&VڌT߳���-ܚ�Rf<�(��Z5�E[$XW���h#	����b���4�Mݹq� α��Wvo���������J�Vo�}�a��"����:)�(��+� Բ��<��XDb�RR�غ?����y��������E�X�1��(�yA����`DĐ3�����D=�Fu���rH�ɮ�)�cO{�0����J#����C����+�,W���4T��Y�a��a�a"m�h�I�7i�����MI������S�K��Bk�#����c/�{�G�|Ӏ�ә4z/���Cx=R�X� ����n!pu�]�����3��J�'6
1)�v�℀{Ԭdn��'/���LtwL�*\m���{g�b�0Q,�  N\��7#5�P���йn�˵�	�w.�}�G��n�m.��D�*�n�A-���՝�v�F16ч��������F��P�ݻ'����ː�,���g��	e�P�g��Ր���@�.�UIk�+���UD��9���x�j[o�}��,�m�,�-]MJ�W�J9���>v�m'.)�A=�G�7�~��U4'���8w��;pCď��c�26�5�Bܮ�. �
 ����h�RC���aT߮�j'/EлWF�|�_�-�.�99�(��Wߠ��.1�	~��Z�:��URB�3@��	I���Jq �!���Bk@�g�Z�p�Y�b/̴�)��_��z�J���	��Ё+���͝~�]��J��±�N![��������CP-��s�]/ K��5��e@k̎YM/ւ�W���?�KϜb�}xLT����|�g�nEC���+���#�D�u��N]�Y�1�k��J|Ɠ�$p=��ްH��ݎ��_� q��4���kd�ټ[��߸��
x�bA��1��*�⌭+��! ����g�/�ļ���Bt���dawV2J���+�|����֞��r�U��Gʡ2,�8���#���Z�
�&���tKH�
!O���G�|׋�Nl��}x�ET<�͖�ͥ�X�"�t����f��觑Җ�6� ��պ�!ZY{eǴE�+�~�su�EY���Ν�������_2�q�0��ы�������-�8�S6�Vc e�_��78��u^{S;j�7H���3�}'�/�ꊡb]!2/N���\���>L8U�?y�]T)�7n�"���hFGk���xꩧ099Y�+++�����+�����׊"
���)��a��vE�ֹ�u]Ҳ���]����V��1��Q>���u��X��n��O���k�[7����0��㭈[������Q�a
���~�$�[)�a@�+�a�QS�S�\�R%3Μ9�o|��j������OJ�;�(����$�3�?�Ww��~z����Q�ǽ����(��i�i۶�]ߍ��a,m�p�D۾�'$Oo*������w�\��_������k8s"���O\�������7!7�J������7��p�����<��s���i��� )�ߵkWaW�k_'�A�yOO��_L�Bi��݂��� ⿵�4(f0��O�oS�6�_�^|?դ��z��:���V�ph���^��Z�R�o�iJc"o�^p��޶F`5�E���W�����آ�����?ceLd���������Y�W�փ|���H��z��>�\p�3���P�V#�8:�2�5JK�P�&{����@������g�ޥ�_��}�ӛ6J(��U����B�����Z���L�0�k_�ȼ�T(
_����c����
�4��b��@���MwJ��<+���Z�;4�.��_Af�-2�,�8g�`��}��0k�)�x��#<��GrR��DN�ʏ̤�cu-4�VV�Gd�eMUUUappp�UB��쿦��X��i	V+r����2�|!B��`E m���E�7��ꢕ��{�Tߍ��3�58��ح��{� ���V&������� .���G�l�b4dQ�,+�I؋���s�ќIg�}���Ʊ�v]�O_酻�_����eE�=���۽�J����!8iA����k���'j\k�Q�W����GM"-�˕�w�(��`��x�b���D)��a:�"�1%���hҢ��}��o2�����ۜ�̈́��v��!�1���AF�� |3{���K��|�wbxx?��ϋ�.z�M7݄G}t��^N��9/4a�i��J
���p���#��?���������(�ńcn��&�K�j	�=��+�D��S����T�n:��00&�d���XNށ&_uY��{�l�J��:�b=.��t���/~�6m¾}��U"&-+2Dg�jM�CYc@ 6=���6�/�Î�1���NEc)�r!jq�}�9��T��	wv���c�Z�g��2��fހ�5˝���lڞ�(fL�p�5߬��v�ک^����:Oz3�b��ly*�j���_���w%s��Ї���T��ճ������W@�7/��&q,}p1��\��p)O�"9C!�ϝi��hRΧ�݆b��Fl���G�-1#CY�|�����z�,c-d
V �����癎�.�j�Р3y`؋�}12\�GD��eq�(������~FciX�ׯ�[�����e�{���k�����<tn,��Pl~+IK�-�?�	����!��q���s��;s�Ϯ�Ϧ�!#�j-o/��h������X�$�x2��ϫ�N �\5�+�\�AQUmNcsIPk�)T�m.>�d�r�5�Ϲ��SiFUm�R�lLE��?��p��x0E	K,T�vK�e��P{��J�-&]w;Bx�r�5�p��H.�31��W���fAǘ������Ύ6l�� 셃�Y�x~�^EDY��lP'|hK���D��%��� �~�X�J�V�K�����c�l�|�7��E��>�����˰�8���lW֬IC����𣧺�ozTy�%���j{i�wo��X ��¥d�tԲ-����=tN���{�2�����۰I9�1	�j�KE��	���`ݖ{V��:l7_��~���1�v�:�rYc��e7JJ�H9ȁ����X�ؾm���'o���3e�"�VX���2a\����l�d���g��h���bM��m+��W���_�]U�ƶ-X��^�D��J��,�2�@��k{E&ZJ���FV汶�ag��������s$�m�H���9����r��S�3����)��S�^��}#J�����'t��� e~v[w��t3�����v�~q��m,�a�u���*�&7����G��a�6v�s�A�dLJ�gfO$��5r�#�Q[�1|��Q�ǐ��H4���p.n��.L�hF�6��k9��_�A��q�V��z�uf�'}��l��,Cs�!Tׯ��U��J���*Fч��	����K�İ*q ��г��܉��v�	E�>]|gGF�R�]�����u�q3�DH�_V��?<�ӣ��5���%m��^բ�����Ѳ�6T�DT�Cj���w��ρ�`������n��n�C1ČH<�s3~�kQ'���k���~ǉF{QE<s��:�1:JC�!�L[���6<��/�C8J�Z�0ǁH9�6	��HH�1�I�K�nͨd��()�<�
�K�5�����w������qZ��}2|//Eױ�_���ɒ�j�'#�:�,k�tw�bk�׫~ȼ��Ϩ�#�4B����y�P���K�tȒ�T	�S�n���Z�����c0��x�+�� =ߴ�:/CX}�'=��f�6������Q$n{y�ReW��d%C�+ѧ	c\j����]u�#�Cs
�?0�̸p��/��I�������)�Stڱ^�ڔ���Ѵ��iTd�Dz�w�It�J��,
E=8����I����x��P{$v��!�tf�^�g7���+�<u]��Gz���Ԇ�T������\.IIO�<x7h��z���aei�<s�Z�m�4�j;��F�h>�*j��⫞6x���£g����p�Qb4����uU�����d��L�E�:e��+�V���5�4~���[[�v�G�#C���Qye�\
���q�#�]l��pU��(9U�l��[>�\�	ܗ��?��e&0��ZV��3�ɖ�g�]T��2b�>�#S�zl�z��9X����8<8����詯V4|&���Q�nQ��$���)e���f�Eo)	�	���`V�s�ҎQɶu��g��4e�K�J�s;zP[Q��>���s��>c,�}\'����-є��V�c]]�c]I��w�b+���)"9�����B[�Nly�bHs�ؚXN��h1�����z��3�\n3�a� h,�
�MH���lҷ]�}p��}\�Pu�H����^p_���~TZ�(US�^���ze.�mya/��Ӝ �b��&nB)�Xt��F��2��c���}tk7+�d;;f����K��*!3�+fX&3���L���oՕ��ѮV����DJh�G4�GM�\ e�3V�
P�t��d9v�U��F��e��Ҕ3kfY�>|�(&ٳ��$jc�����L@�j��j���Ud
u(q$�5�
��9�8�؈C��5���^6qX�6�#A��W�/L��?ލ���ׇ�C?F���PQY�A�&b�=���O�P�@g�&��u��A�`�c����^���Ub
�zϟ�"M��[&�1\|�4^�Ԡsb �������y�^\9�*�Nx��g����X��e~=�F8�*]��(Mb����uXj�f'�^���;���6M�:�άNrj3�W�}�S$c��{G��g�zE�8�%�S8w�I_#>�;���O��Z�!��8.3���Eh?/��Hʆ��l��H��k9�9��DʬĒfMh���ݝ��
|�f\�k�St e p�]�RH�P�B6�B����ԗ���x��uY�F��+�`�W�\$�Ơ/�~oH۳o���"3������c���r���n��}U6���T���Pq�u���63�1�)�YՀ$��r�/R��n����F���
b
��}����3E�w����=���=������Ug��f�>V�)z;�}�]�����	q�Ãz[F�;����AUU��`�WOS^��~1C��ߢ���˽�a��mӰcF����������W��']>tt�@]�1{��!��ߋ�	F%����2�D�Q4&,���}����9�~�Lѻ 8	�=��s��{{���p/ܵ�b1z�.c�w�����jf��\NkKb��Ӌ�7<������ΟT�v��qo|C)��"������	�	7�g-����1�f�C�2�"�0��F�6u���Wr��Q�}����U� v��%�����^"\WV�"����$.U޺cf[�n��Mݲ�[$F�P���I��]��.�O�]%����G�/���V�b-ҊbY4f�c�L�m��Ռ���H��ַc�소���5w*4�r*��c��]Uׁ�5۰�wR�Q���Z�pմ���� =��
���*�	�%&T(���dW�)z�_{�����}��)�'|2I��[G�[w�D(�h�EHj5P�:����*��jE���\ e�����f: �t����V�d��W�u�&��ʠ���k�kYJ���},�)��?:~Q�x�R��p�O�Q�J�^H�-
ӛ����Ci;<��о�X,VI�phP���D"_����Vua2���X';~)��3���P�<��K� Lgr��r^�o��
oڌ����o�)�Ks������3R�5H�ݨ�'�Q~�5to�55�i�-�}g0pi�lJ�D�ָC��mM�:ᙖ�I��1CK0��A|า:��GtZZ���Xچ��8ۀ��(uh{{��I\<���{�?�2H�\z�߀ϞQ�\u�h�����˾R�:5hu1��YlM	G�Ɋ�E�Kuf0ӧ?Ňi,��,"S0�H�J��U�d_ĉ:s
�S/"0q	�V�;a�wx|O������^~p0Z!%�7G�hzC+&�b�z�"u�,b�u��Ŋ���|����)�=��� WY}M=��}QN+1Nѭ���l�N���A�@��|T�DZ10�3B'��Ja<k���-�Jʋ-+;h4i9�w���ae�>���y4z��s�11���t�A���e�(����U�<������Y}y��Kv����`�C��FUV��"ӽ}E�}B��E�ď�fdS�w�s3�j攼�c���!leЙ���7�!��U�f)��a�^h=��lX҆Zx(&d�7���|(��3c�b��+�G� P=�ݸ���  n(�������;�[��MӢ�������Tb�r��ʔ����J���0J�9!���!�'c]Zc�=�ϻ��U[����ط"�Ğ��x���K�ja���#���mqUH�;�}ؘ�Bf��/�z��dZ�~��\�נ��S����=��z�׀����l��W3�m؉��?���Bo�:����2Y��Oy�̷��mkĢ f"+�2`�ޒ����)+eFn����D���{�Cx��Ö���kg��l�����x�e��x����h�ޣ�Tg}�0�"(Ґؒ�Ծ��8n��	e���oym�l�@~����bʏ>xLY!3���o�*@��xR@A�����	���s�b�.�b�"d-J��ݬ$� n
��3��۔Ψi��٦�s�hn`U۴���i&��O=��-u�R�I�Bk���W����R>@L)2�^Ō���3�K[�X���D�͊ku�j�z���[��^Bܖ��ʎ��.�RLE�eD�ԇ5ϓ��+�u�w�m�h/�_V1�����1�*���a�\H&���{�}�M�s���܃�z��J��^�@;7W�FÅ���
x���$3�
@ʝM��7��wL���P���D{g�
S��L�r��KW;�����n� �$�g�
j�Mu|a�2ū��-s��+l����'�ҾY��ӆ>߄ )��g5 e�o�Z�"�X[�����T�o��f至��̠� �:�J�d�Ʉ-W�UӅچvT:5h�|΀��s�?����⹊�����j��c?C$8! �&�YjPG.��#�a�nՊ��=}E�M�sc>�2�=�	�_Ly����s���E�|����qSG��rz�'�B�u��߇�c��ҹ2�>�\9��}v�N�ϭ����@�rT��5�����$�S/Ë�VD������.��o�=�]o�\f胢�m	��5ؼd5͌�����&�5�&*�F�N'���Q7�F\�#9�J�Ͱ��N٬�����������h�J��bJ^K\_f��Qס�F��Y4g���xY�n����Wy�y
g�N��^\  ���Xm����y혱����9�T,��~E@��;H�j1�:3c���� �l^�y�㑿>u��k͔9̸~(z}�NI��`) e������4�Ld삊Q
}��Ҷ�˯.Nֵb���2�̔�[u�x!��@�z͆,�Q��]�?����4�\u�[t(�Ao`�q.>��A�V�����c��^�r��KpS���|c� 3z�Q<\9�.W)\�	�x��8����&�xF�!�d�<��oh�Ɔ]�D��^�v��ϼ��3���Vi�b�Hn�F��C�־�Ɠ<�\'fX��y��fIK\�q|x�m�%��Al\�k�܋{��;����Qz�"��i+��Y,���̇�UVl��s��V�5��;>�t2�{��V��ɔPC'��!+��w�I�*x��u�������$�:���R��n Ʋ����a�[>���l�����'���R���F4�-���z�zz[4�c��u;en�Bْ��E���5h�]����1����+����7K���d�O�� �!S�
+e1�\g�a�}Qr�X��ڥT WHc�N-��� Rv���ܱ�_�[�*�ܬ�|�p�j9U����p��  ���[L��R9>4�-M��%����u��]�)י���\���A�I�@k�)��IH;�z:�k�^�0�(��A�E0�Pp�h�d��Q����2��M��>�c��pT�Ο��#� �|\7p̅��~XSm�_4!�V^���!�0!��#�@MC�\�(�#�5
�r��k�L�R�5&'v��T_�o�a�D"���p)nC Ch�,܎������H���1�ܯ���=5[��i+@ʷL)S����4m	�\ӸN�[S�Q���p�1�G�<(�@S�`̉��l�A��{�j*����/��P��l��|Ѹ��L��2|F;��^�)j�����-�]w?������!��kCO��|(Ë�Zt��`�����,?%���g_�O�b�s��Y����Y9���~�r����h �C<�Wr���j�ӓ�K��c ��x߰|ɔ�ĝ�ȗ;�;�"i�-�C�ۗ����4$�Pʆoy[�k��]8�"�B���mx6�,�7���$�e��e���≩�0�q�7�@,k@sIF�����D?��쉬p�o��7:#��a�ro��h�ڬZ�e)}1�n�BkmK�����<��^:�l`U�'�e0?@"����4�>�yL�D9�L�^�D�5�?Ĝ_Ӿ�_�1U���h/����A_�Zl�'g�Oۛ���lnVG3�]=�i5FV�$��U������w�h�9����^=|C�q�)+���ņ�-�,�d
��\ح��.�zx��\�T~v�Y�1@���Jv�R~�Ý{�񦲹U	����aS��ɀ�Ю���_�Y��ϸ��2Y����������4|B��.SJ�Ɍ���5o�PJ���
�8|������R<+��@�,��̠i�Ж5bY�y��Y���c
I#����o�gv�`\9��D��"h6��c�ϟ�'G<�_r���7H�ڲR<����?E�]e)��=�����¿��ݲ��~�Ox����n�G���l>K��cI���	�yT��Ns�W�csi.G�L�qe8�v�Hu�wCx�5�{�S��t�rd���!�:i?����uO�Xb���o���������.�޽Hp1���R�Yf�"K-f1_8{��_�=i8p�r�t�a�����A�L��g�T^r3���}�������g�c��~z�����=x����qebS�2y���t	���s;�_��Ƕ7�n}��&���;��c/�=4"!x]�C�Й۝1l��WP���e(B��^��JW^��MN���F9�;�<�k��.�8tfI�K����V����}xt�Z����⿾�_v��$�'���Aʵ��:��C��b��f�6�Lf�y�"�y�W��uRA��}�y�w�n� ��}�L.yø�9�͵e�q�a�W�5�7����W��A�WNE{9	����Բ5��;J*e!��	�۱�vl�>^g5�ey3LPj��1����YN4��M]�Pb�[����[wsG�݊\!,I��O���Z�+�O�{{�%w�
C��t4�5�O��m�2�o��"���:��^EO�N\���cS�;�3���XB뚏�TMl��+a(��:�5��މ���q<�!����-�p5ʇ����YlMX�,W��e?�@�(������K�{��7�yÄ�����E\ڄ('����ch@Z���b3��x!mWh�� �x<���ާ��-������T�g�WW�Gz�0����_Zp�P1�	J1L����58uɇr%��uT$]u�0V��a���ڒ'R�T*,�I�Y�=���˙�LƑfy��2)nnh����]yp��y��V��iI�۲%���q0`;�i!G���t�L��@�N;�%%L�@��@���f:@&!)�6q�����6�2�й��]+�n����Z����dO�̼��c�����}��}^�H�t��}�,Pm$o~E��%�����*���7�:��^������"H}�]�{��Ú-�<�3�㟞8�}�5���3"��x}��.���n!ru�-��?�S��M�zev�M/�a��k�%j�]8ٺї����Z�i��NV*���Bw�����,�~�v�,�O�[�C����rh�a�������B�V���(�-�<f�&���/�w1BbS[U���a%n}g�(@��e���4ʗ�ӠE ���\��|���B���^v�6"���Q�����+�}>\�{M'ph��~��+�\*��y���[�������b�EJ1�:����,�,ǉ+�
���^β3�Ch��&��ơʾ��*@�r�#r��>8�k�Z�99y�ۑ�a4|�&���B��3C�N�b�9�bܭ8Ϡ[4�j�:�v��݆���p�_�5ř�rn*����ht��f�+6W�bIp]�>�,������g�:<&06A� �ٽ�v�#J�����ӱ���wM�8�Q�U"��xZ��y7�=�l��5܅~{&��\�\�W���#8�Q���B5zcg�ZW�s�z�_��{:���:ԋ6�����;��{���7���w �r�+X��/�`�E�PN0�߆Q�Y��WcLQ�^��Jۧ�Vb�� Vt�W#�s"'G��8�����]����F�����VWh}��m���aDb$#H h\$���AW���i�Є=jq���)�z9zO&k}F��L��v��|ۤ�Π�#�$8ۤ��	vr3�6�)8+g���L�Sv�o�r�U�2��͡B\�R��u�[��}981�R�턅�iο1\,+oeD�"�D��j"<��ن�r�<9.Z�U�HR󍩬�T�9�G8q4��f�>4�S$��b�G�wR���:�o�9��n���q�L4�����H搴�F���H��#GT7�}V �@���k�d
�����Ao�\zT��TK��u�E������T���M��x�����M�[�'UO���Z)��#�S���s~�(�4�>�ͮ�l\6��.�i8�ܨF�9&��=��Ry!5Ւ�Z�=%=^� �)����י�"\���o���<:Yg�>�s���W{���*�2��8�Ӫ2�h?���oFIf���Z��}���`��E��qP5���A,Ms@�a��{0*�(O����E_?nط;�l���-�e��&����kIi�=���"�o�B�G���xщCf�r@���R�0��FM����AeƘ�8��;>����p��k�sE.�D'#
;�{/�\�I�f�%�ıX`wd਌�sԡ&d?�Q(Hs�\��ъlȹ2�jeВ6~��=K�C�}�Eؾs'��b+���L�R���̬l�9�Q,�� ��L�/*4��
��.�2kw� vd��(ï���q�x���x�ָ*w �����kP�|c��F3�\<�U�#�i��\�1nپ6윫))��E�Ox�v���!-��x�	��L�b�֭ؾ}���s ����&��1�q��������yΌ�ЫLی��P5��B7��F��f�ʬ!��Ƕ��nkYی���Q|��[�]����Z�Ҫ�B�M�~�>1�����|����-M������S�`�`�ħ��f�o�EŒ���]�|2z����>��]}ʖֆ���t5o���՚}Y�Kk|����k�j1�G�N0�WqVo��_�1o!|"4��Ng
Y�I�/�.����l$�b4��EK�'�#��k�u�:s��.mt.�Z[S�]�b�,�^Zc�cT��n�YZ�k�]��D��u��/�J]��)��ʠL]'�6'g���f�/-<#��k�n�P��-h��ҌI�2����1� 7�5���ԍ�Y��yvfi5C	 3�6��KFF7��[V�d�²g��Tx��E �eɣa��'1���/n��ӷ݈o���ۚ�:e�-�sm�ǓV�5���Bog�R&�2���NR��v7�w̯ˤ�b���sZ�@�9��U�A�� �%!�3�m���|��'�H�Bn�DB�Dӻ��5P�(3����6��5�*���׭�ҍ��p��24v��V/2c��Ԭ* ^�w�\�ϾHo/z��5:��_wT��n��WX���v�7���Q��z{�ƾg���1��=q�=��Cݓ�B��r��p%� CCC8r��H_h���뮻�m䄑d �� ��7(#���L��*���m�H�� 5B�$�
^��O�ѵ�WlVe����4�?�����IT���������w�Wym����'�۞4+AYn����~]���z����Z���mx������ۃ�JY!{r��46����e��|�ǲ����-����5!#X�k6W���{��U{Y�������D��!x�%t]D~Q��Ɓ���������ٱ��oʏ;'3p���M��K�;aӍs�����ܰ�
?<|R�X�0˩��(��%PQi4Ӊ�0QD�����0�XH0�y�����ڼFӔ ���s(�3j�KOl<׻����[W�Ye�n������fx{y���\݄�SqDL|_��o��sǽ�n�6��Ki�R����*锠�	뤪��>�X� ��6�+��fK�E 9.�z���;�ke�it[�_`��.Բ��i~=��HlRo���r��ru����=��[�7�0�m��|h8�`��H ������2��<I��^�����XV&�J �/�z�E��[�S؍g$a
3)a���H���'�/�s5��ʤ�� ^��!a�]���"��V��
T� �#�z���% ��Du��F�d�&qQW6�K�{�E�₨y:[��3�����B0�z�!�P��� �^FPÞq�k�c[�Pf�
)7�rpz�`Fɒi��j�n-lEma��V��æ�-]㥁2�X���R�}�zT��i���n8E5d�U���3����`6]c����|Q��������VC��G������.���d�>���gݍx��MbrLS{��}RKkl_�v܄�lk�h@L��~���j!3�"���t�_W����;���z����m��ΡT�N�[�@}bX����K�l��:�^��vj�O����!8N��tUn*�C�w`wv֔`��k�������r�U���3ޓ��h�Kg.���R����7C�k�a
It��縃A�	)�Iy�TS�d"Y3��ŀٟۅ+6�f�^���
!B�:��|=������W�{�9aK}�se�v�����`����%�NTTo���C�}=��A�DL����74-�0��Αe����֖�x�=SVV6g�6���������؍�(��`�s�U����>�A���YT,�6��_M�,MG��cˑ.1Y\�l�Ṕ[��O���ە =�Q��z��&պX�YB�ܱc����̍R����?����9�R��"��7��kBc�I�P��|��Չ̴����)�A-�^܁�63�W�HY�7�v2շheR&03�������q�2;�/�\��9s=�DH%�����i$>�cP 3eܖ�p;�V�V�L�-���nF�d�&�O���Jw=�ZΣ��YY��0��wF�����Hvh]\@�Y�s�F�.����R�Ő!LP�%qg��9m�����aY\7��e���E���安"�!ZVk��85Z���2���� ���E��d:���A�#8�хׇ��!хr�z�?�/�r���J�BP�D���k�T��L�����.J���qR���P	V:��v�'��݃��%mm�������[2��)�}�'{���:�d�م�fp���/��]��ﵩ������d�7j\�L� _�J
����Qcb��3�lj���9�<&ˊ�l��T�l2@A����̜��4Y�6`������I�YK�]Q���Ƣ<�ٿ�T��N��_�J��4���������a� t���/Kq�[�2.���;Y��#<���{�~�ӛ0>a�y��Td;�� +\DxAD�Ud���M�R0����ĉ*�w�ܩ�&2��=�v�
�6��� VMM���oM�y� >�����ǯ����:|���زe**� �566��߰aCX{��*ǁ}�9q�]�c���*��[dG$>~*�C��N8��e�S.�&�;�f�G򔘅�i��O:�ʋO�G����ÿ�g�j��OW���E��*�(
%�Ya���>��F�~�i��W��v���Q��3Ϡ��ZG/�O$S�]�jՌ٣�a�����E�����+���{�w�y�>����s����#�<&��3+K�9�
a�3ٰ�<|���^�||8�5�}?`Ǆ��,�>R/��5<������9b���3!(3ΰ�HDr�e��8Z��y��D��bB`Xg����oy-���<�\���^��Au���Α���$\�4����	`#�KKK��k��"	����=/��,�/.AX�Y]eX ��&��`TY�611!p�� $�\�9>9�;�Qc)�uC,D�F�w���E�ji_���ٳ��`�'#�˄	ΐO��g�<#�Ҙ�E�o����E�M��J�S`�8#�/�} �I\"0�^*�====J�� Fsf���ҫ�B���_2'#	B�ub�f&�Է<%�Fi7�G�2��U�q�'�v�?���%��A[HY��#J\��4f�S4L#�+�:ǐ�L�0������o�|�D�قU�`\g		���$��\	b�?��Y���c��O���Q>V�vg7e
q'�G�c��Ĉ��k��i���\\� Dp*�=409�LZ�%�f�7����ރ��@o4DD���y�������+i᧕�G�q�'�C�K΢&Z��O��!̖���AZ�-����px}�}#�]�h�z9�YI'��MZ*��\��1�O�����>ĭ�aB�FsI�U���7<����yi���j!M���u*��E6w���ۤ� �E�Q�e�|�9�V{�!����4Ї"��%p�����1���)0�4�=%��+H�Hgc<0�ԜU���(���Xn�q��v��r�$@�='���H~�+�lND"�'��#o�e~E�-���{�X���؈(q-cL�]��^��Ƅ|��n�M�6�3��X(��+���3����E?��W[[���v�]�vzDOڐШe<�Dc}���oN�(��c��N0� �`�s-,v5�Dx�v���<�܍�[Y�!�hd���y�*q�1G�ƍ��SO���qMΐhGd,0���&Hy?�����~;n������}��:��t�k�g�)-C��M��
��$+fG|~W�s�?�2�"](��D�K��"�"'A��TҀ�}�QC��^Þ={�nݺ0q�	�o)�r~$}��n���ٌ����a����@��ov>�i��'&�ym�jݸΖW_}5&["AȊ�ĸ�٢�]]]��r���+�����L�;v�y6+=��|����('7mX�����Hnmm����!rA�DC5�j,^knn��Ç5J/�n��__�L�M���xg@��|����/��X����=p� �x�pNs/y5��"�Sq��]���E ;�]�w�x��򗿜�pT#4=���g��-W��x����g?�H��U�b�_ ��y~~~~R�׬ĺ�k4Vnf �tP�Z�f��p�'J7����� ��rd߾}ػw�a$�wܡ�Rq����~���l�-�ܢ-:�$\���j�����&OG���O����p�f�\"���/3�J�Kau�e ����$�]�,�^���*�,2H��o]��.���)�xH�X>��]�f�*E�P16�X���C޿"    IEND�B`�PK   T��ZFǫ�>  >  /   images/3db32f6d-ca85-42a8-bb1f-49cf601f6ec4.png>���PNG

   IHDR   d   K   �"�   	pHYs  �  ��+  =�IDATx���g�e���tﹹs����$I A0�XP\��鵬��6]��Z��\��$�P�T[��k���b�MrwAb�"H� �{z�{z:w�|�Iz����}�1�+��Ew���7>o��c�_}�ڛ������l��˛h5#���80��i �����ض��"3���յl�ee��`f���oXN�cۛ�m7�^�
k�|�EV�P,n���G�k����1��{ �߆;8�oQ~
na<v6�n�CD��r8@˲���V��0��<�ӱ9N���P���A$�yz�a@�S������}^�r�<���a�Y�����v�E�~�H���,�׌�^_nb���/�A!7��B�/�l�D�P��W@}�{,ʔr!B�D�D�p�d@d�cB�$?������V��N�p�,��wt� S�����5�(��<۲x�ٵ,��d�F���W�/���o}�X���e��&o��Z9~�����#�B
F��ϟ�'1��L�j�;]>3�1���oَ��y���4���A�QL3_�!��f</2-�p�M�x�Ї��$�L!)�Y�roȓ�CY%���qpQ����tm��G��� �.�!�
�kE��/R�M���H�^�;�*�����s�=�mtGM\��$C3�k5,J`�0 |t���M.�/���.�6�(�G{�Z�>+�|e�(��F&���s�0PHU��g��jIC�pG�� ت�͆�R(��n�Us77�)�%�_�;�͎0��s����IN%[l@�&�K$<�:��x�X>�H"��l6u��+9�@N�d������g���1UX���X� ^�4�`���#�_�������P�;X\\C��@�j��P��H��Lå��pi�#�E8�n���|��,�Z)됸4Y���J9�R�B�` kS�B!<��\�������k�/#�R��W�4�i�@E13=����(R_.��ܰx	kی��a~�U
[b��	q�5g"̶�&>O�%��fj(?D��m��6���D�
��,�&P���G��E����	����mu:����
�V+�&&&�7Сdup����.�G13��_B��`��D)+�u`�>��\���ʃ.
9�����'�xS��(P������P�H���9p#[�3|a�:a�%�'�<y@����?��VJ}_������� ����m&)�3N�C���*��k�����<�1z�0e>e� G��-�j���?��<��V��w�`o��#����J���F��<\zo'��TG,Z�Ǳ�3hu��'����4H� �۱<�7}\_��ּ�5��I�X��hwC:��ĹYQ[��
P��f2���e�h���::�hڛ��(�.���mJ6�'&��S��*q�e��O5��8ܘ�F�Y��L����]4.ٝ0*�E�b��3S_3����U+L���5S�����8�3�N��dqyv6��/~�k^�7�IH�g<,��}�vt����,2V�C��,�\�>�Kph�����MԮ7�w���$2���+�1��ں�����N��b`�c�e�c�_�BH"�M�i���K�&��&�-����q�Il�ߪ�p�<6�&Q�Ddt���'E6����0�m"���/�cm�c��T��3f�hk���?��J/�P[��z��XC~��_�Yk�.�WVp��������������l7g�h��|.�-�P��6����Y]:�so-au~~������ Za�]�q��U��ֆ�0�_D��[���p���(Wr4m��-qjt��H��.�Y]�����U��M""�4�~*��[��R1�b����.1�d�N9�l��T��&���^m�
Ko��|Q�(��13��=�������ѣx�����;o�Z��Z�����o��`��<�?����+��=�z��4ڶ�<��8�gat��ܡ$V����iu۴�4%$�x�p1�B�S[���<���h�uiV,j�Mo��s���1�r,�R��(?���7I�#dPV��DGJ�0!B*�1B�q��s�&��C0�CD������\8N�q�(���	2�Gb!�]�°$�0֘�ُ�.���+�����37������.��gHbZ�����<עN���ݵ 5B��x��!X�:6B�=����Ubd
]X%�/��r'�P[�E#}�4SEJ���\n�N�&��O���Lb����w��a�3�)���	�X��	�	�ː=m���a��≯8�3�8�=Հ1�Gk���-���n��S��\Z��c�qc��IB�����@)��BJ���K�k!�[@�N�2Id�����dWP�4�+�o�P�)%A�`�ڼ`$�$�V1O�$�uȘ��0`3�@6?LG�*�2T��|KQV��F`�X?4�x1FS��1RI���VB���c�w��>�2�ה�c��>��_.���H4���084���������r���<l��)he�Ƶ�F8(d�)��#:Z^0oc|��f`�U3����g�}	g�{����Pڻ�)T�i�2-[,�ۋ�����`�P�	T�(�ԯ�V<��O��J�'$ԎM��!"��v�f�#қB��m�ߕ'�W���0�ܻ`q�-6�+�H�RFW�S�ݨ7����_�K?�)���k�,P3��4I.#FN�FK*.�R&$^��'v�1�7n:<6��G�jMB���
c'�Ӟ��̵UR���X�.��yd�%hI����Kd��E$1A�-Ͻ�7ػ�!�bX�_��Ð���- �n�G299�f���188xsuuU�����6��G�S+:^���M�v��Q�&�A��H$� ���L1�l?�>�d��m��A*ՊP]�0$j�_9�2.���Bp �C��\��Ŕĥ��ˢf�Լ��ky��U
�G"����pg�Q�����>�Cc��A>"4�K�����ߏ���Ŀ���;��O�����j��VI43ӎ�=2t�yjC9�B1׊�oj��ӟDF�˛�;��h��(���$!�8�\᪷�D�"�*��P��7�5�>ɠ �0�p�h��x��q�&k�f܎1���s>���'��
,neH�=�bQ��}���_	���?�<��s��C��^mP��=�C�Φ����ɹ�t��U�ބ��� �N8+Q���+%4�;�Ԍ��% ?R��ѩ]'j��$�A�>�Qt؎�� Ҹ"�s7%� AT�Em�V�� �����AnG�ߕ�wBq��-�B��Vj����׾�5���?�c�g��?��ѣ�Wa���i6�;80E$$�d@	9O�W@8���t�y3���]:�JC�^K������w�h��{
������A@5	��I#�؁�1�;�Ƞ&�KDD��z$#����e\w����s�`�ۻm�OK����X�5q������`Cc�sm2�~�ӆ�+a�Vg����F��_t���Ѧ��W\��n���h� 'M�;��k��ׁ��ظ@��I8�v���D�/fJR�k#3�,�xx	�-22.��j���3Խ�g7�RF�IP�I?���q��m�4��k��y�666���>��ϣZ��cٺ��0��4u�{�����a3�Q�v~a��#{Ld��"�m�Z��q���O���Fs�����uޅ�CI'CL�͞H���N o�I=3��𜜢8SAE�yM���v�{'i���c��?	#�t��c؝ ڒ<�!���c�$d����������Ui���y�hjb"������ܨ�4S�Q�q18���{3hn���s��-�.n�	Vi���q���M�]u�q�!�BrW6	'�$��U�S�3-ήj	����K��>�㈼��;�����?"1ũ��E�5ڡ�_119��]�(�>Volaz|�f6-�=���|��>Xã�M�����pml�U�-�����B�v'y��[�&�,�*���D��gD��,�i�h;Cj�y��|��J�UaR7���?����n	�v��}���ľ]����(�k����o�Z�ج{��x�b���U)�M,�l�r3h0�_P���=�r�(�(y���j?n�����[(Ь9<����ז�Z�t�Ȕ(��M#��hk�D鄸0$'�X�調�M��Q �4�������%����Ȥ[n'���F��ݣ$es�?����ws�s��M|oc[��]�u�[�!���z���	*#�k�WH�5�� ڮ�IH�-���F�\Fa����MI���kx�a����q�w͎�V�rߥ	*GG=�=�1�8a�ŭ$G���*1��$9|ļI��Қ�w�����d��ô��߱yI�����xi2.1ʾ4���|�:FRJ�a
��Lb��h8�`�����0Ē(�k������ݠY����\� ��K�XG!���͠���@i�m��dT��ب�"�]���)���鑁HA���$�Є
q�g��K���	�C�k+Ӎ�$)�z���uW�\��hIyssS�I��g�Y���+biӼV�U��Jۏ�{�p�P,auu�?� ���#�����W����F��d�mwP.�z��'O��"ו���u�]8��M "|i&8I�[t跨�ݪ�KO���0E�`�q����F"_��y��;h���r�'hV2ȋ�*�������bu�N&���v
ST7�E�8f��`�8}��:8|��kW����C�T;���M����x��G������$��I���x��3L}�����ܜF��z���K_�"�ޫ�_~#�c�ڪQ|4ȴ���>� Μ9��y�&�|�M�:u
sW���ٳ��K�I?1����~��
M��Vz�Ξ=�3��v�%�hl�Fڅ����q-;����9��� �g�������Q$���5 �
 ptks��� �k���B"��q�D�A��X�p
�&}�y4+�l
�%վE�%-D�VVs^�z3�#ǃ�>�/R�~�aJ��������SԒ�3��|mA
5ay��Yllm�^obue������E���o���ޯ�� Ӫx�ש�6N�<7-�1=��Uj�>��g�������G���+�|�2鴖R��!	�H[-�5l7nY���:�P�@`�?�k�~'Ծ+�bM�tx��c���;!#�g�AH�v�`����*�6��=���]_ǉFxN@FK?A"�2F�	�_�H~6����E�R�4���9�-<���=zD5b}}�����
X#������Z�&������"���;�w�}ǏߍÇ�`yy%���wҐ�a�G������?��D������&�Z���K�	�x�y���\z�*5�������7!qGv��2��YG\��y���E��aπA�K��4��N�;#�%��?i�?�~$��O[<_�U�[������kah4�W  �@_�y�S(�h�Z��M5/�y�:5�usDx�ԧH�tppH�-��x������Ьͪo��X\\Tf�ٳGm�ԹEK$@믔5���[��Ć�g_j��'��������+/�F�<FsZ�5-�ۉ�S0L�,C��f�>� ^~-��'�&h-C"%S$�d	<4���m����ϣh����2��ïyZo5|=.���r��B[�h�Կ�}�y�V�ė�bx4�o~ނ�tp��tI��y���믿���x�y���J���O~W�\QMy��Y�~�������3q.�E���oR{뾧�z��[H <55�1���3��¸�8Њ{�E��6��O��d�L	�/@�#nE����X�sK�b,�؆���z��\yo�����UB����Dq�!�R-�m���5
0�D{�ED�?�؈�!-��D�NŁH'b6���jC�3$"�:��L8@��)>��ӿ��ݏ��זB�[%����o��,�969��%Zz��a-�~�+�P�x��5,��'�S?!�A��O>A�UP"�۷O[���s7*��b�����1���q��A>���@|��¼4 �'?�)&�a�~\�|��{��	u1R��X(�vP-����:���h�R��i�U�Ŕk�8�|��/�{��/�̾�s�bs}#ACD;�eZG��L��r>���M�X��H��}uI�,�f3"|�O��%�<��X@�S��4Yy
���vO=3FIm��~�c�s]<R�bӿ�����h������H�:�}���*����<p�����/��c�D<}��j� Av�Ⱥ^[%�^��_���X��I���߾�6�^mh��T�> L�v#�o�x�}XY������I�6�=�͈TOĒ��@��}�?�}*�/���wb��nF=� {��ی|kq���{�������������׻�G���C(�m^XT�Z��1��6խ�:X^�c����H��~�SS���a���G���{sT���Ьy��g�1{�K��F�+�� R�3%J���6I��$���}��6O;}.]�L�3P,��-|p��J���s��%����XҤ���_�/Z�����B�3H����K���y��'EZN�Z���ܹ���}-�5Az.�~�b�97S���M�U�/\��C��m4n��j͡E�m��9�?�gK�~�x�Ց��<Z��A�����F�Q{v�������2�}s�ji`�?K���k�DX���0NJ�U�m+��Y��*�r17[Í����++s��X��"�1�?kd���_{������� ��N��i�f[�'�%;y���o �|��F��YU�ͺ��Ν���v;ǿc!z����)���B�����
��מ���A�Ih�Esח�����vUS����b*o�Xb0�)5��Bִ��Y4��"��!���Df����I�P�&%&53���;(��>^�{�-��-�3��������$#ejT�7��	4m+�������*���l�11IDd6�u�d�ܟ�`�+k���~��D�$��Ym}PiL�t��I%���,�`��,�G5J�H�{i���y��y"�31Y]Q	�\�5�z��WV�9��U�h�ν��z��J���ɪ��juK{�d<���؏�8�=V�9M���k�jV��۬M�eҧ8",�9u���{��<ͷvcF�Z�ڥ&T����}4	�F����1��gx�t	e������|h�ii	�C��I�OpwW�脧Iµ5�ߩibu�AI�0:���hR*x��Ob����]���W��Y��:�����za�j�!�D\ׯ��!F������/��Ci�&!�>�L#q��Je�C߻wL�z��R��H�cD��V�73��f-� )h�d;�i�����4�y��y�7U��ܖ��ި5~��Cο����+YS����r���u2�abz��X�������+kulե��Һ֥��گEkK���z{�@1��D��C�o�Щn-3�l�3��?`PȀ��u�5J}����!�0���$��ؤ��hꪨ����#j�����>"��/Q�g�4���H�z�f=x��"0!������.�f(ـ�>!hN|��C3jb����;=��g߾�$�{`�N���xMo�]����J��+I�nQP�[|H�v�ح�n`bd4O�t��:0�N�5C'������:��׏�s�؟C�f�8P��(���"�}9�89�>���1����0�%ڿ<�zw�UO}���(Yv׮uA�N���|G��7/���}o��j�FF��7/S�g콪��k�R�T�W1������e�a-����2w�G��$��	I���q�� I���
���@�ݙ���&]�'G3>���3D:�;5��.L;�ϻ�H���Q���ކE�g����k�],7fItG�$��|���ΐX����7�JU�����Ξ�v���Rc��,PB�a��E�������vS�������3<���Mm��勵�jB���?K�V�`06=ML�&�J�W�/�.�C�ZR)��6v�W��Ro���M�.zi�]2�����Q"�+
�O�<�(�5Iq�\.o)�f� ��X� 0`3�lQ������mLZ\Y\04R�䘃�����Ɖ���_\�� #}B�-r��G�.������8�rND�Z��c<@t�7u�<��סCm1��״��U��|p�]�}���|er�ٳ�i�Z
1oܸ��� ܁-��)-��m�?>.G���;L�M1���%�)�WiR��o�4=��D�x���{�x��)D;z�R���ʐ(����#�@��k-m��Y��|B�����t�sU�蹌�˴��c����`����遳��6F�u��Ծ^:�1�	f��`�����Ah������� ���j����<�WgM?�'�/�J�_��Up��:V����+���g��v�D�yr+Q{q��(��c�vǉ�w߽��Q���qa��p�..����L�h/+5������w�Ky4Lj���dX��z��)/qF���Z�m|����[�����[�u��� 8x�E�������n��F���0�@"ָN*m=A'������ػX�c��D�f�Z�7P��mM����ٳOϿ뮣N�(����C��V���06�`Լ\Z9��L(�}�e���|Tg�n��S��u�{�MQ��~�����G;�/Ԏ����)��H�ڴ�O=�y{�DLǳ:�t}��/<��n\����>�����k�O��٠c^�°2�ӥ%F�^'Jl�������(�]��.�.9�{X.�Dm��S����Ӕ�������6��-:xǏW�������U��Y��f^��Ęf4��xR�$��>E;c���r;�����0�w��q}=V�[K�t�q�R���ݵ\�����f��A"�n�8~� ������c�F��������,\
5J^d��jmh����<6��N�<2�=�;� ����+m�4���^���gGp��*������2Q��2���9|��G������ͭL1�/5�cǎ�ܛ�0��οx*Z�%�r�^���cZ:�H~ʢI����wt%
I�K@�JgL�;��~���k�HgZɭ��f	JR?bGflo�9�_D�7��Y �^���=x�g`��F�$��3�P�.F����,�l+������){�A_��k�#L'���&�`����&���0��1I7��#wi����>v��`�aOK���D$H��A��w�yOk"��~�!�KR�J$���@��/J�nܞ$_���6�~���O���j�m2�����F�g"�P?*����F�����Al\Z����/�%�y!�s3Ԑ.'�C�h�}�"��!Y�P[{��]���.��#�Ǖ�[���L���iry��-b����R�lUi�j���ә�W�0Z/����=q�fe��7u���?�5Ik��I&J5G*)�Ç������Y;&*����5cw�)�m�v��%4Y1Y��S���Eͭ*��y�f'��HK�:�}��2��97h�,M�u��RmO�+��ߧ35�lR�utʂd+,+nK��� 2�AL��6�W�4Z�.!?h�ku�7d`�^�\Ѕ+�БCx���P�ZW��-5O�"ձ��ˀq/���&H�)WJ|]�����8s�a��6{�
F�G��R��B58ط��R��H,
o������0�n�=������=��^��nL�R(g�V�t�]`s#�����_�9�Z�g10jcu+T�?AH\'W�
��化X��}7�L���J���&Y�����=���b_��8x��(;��ѐ�P���3�L��ڣKm�ѴB྾!%���T�9����ۯ�m(�*�:����dt� &krrc�<��qI�w�-5S2VA]B��e����HK����X��t�(�&D�S�d�؏b��t���F�d��D��ʐ���C�,H�,�D��Dmdy)����������L#Ğ�]��+�ȌJ�m�/Γ�Ų��JFdiRl�'߇��dt2ԅ ^��*������*�&�5(_���������u�,�����F�����x���|��{������V���q��U�<ysWgՔ����g$���
�WO>�5���M�{�g�a�8}���v�������O=��~�:|Hc��&$�ӷB�ݚ �L!~;i��ѢZ%�+��O'�i�#��72�5��8:�Q�\[�a�p9U%Y�����N����&29c#�:𛌘�}�.�Wij��8�$��t�Y��X"��F��$�;o��һ�.j��F���:o}�Z�Km��Ik�t�CC#8s�Ο� �N��1u%x�\�4��#�ui~)��5�:11����$}���R����՟��s8��{�W��ѻ^7���RM��:YiB�Ì�����A���m�}YI��v�ݪ�>�A���&g|���G����ӶW\XJ;Q��d�fX�x�F����RM�R�]Y&��J�{۲�U�hQ+�e-� #�2K�ۭ:N=���H�B�����V�<o��{4i��T,�W�=S��}�;�k����?�����j�Wʫ2�[�H���߹���ʕY������{�k
u�����__�B-{�cAU�%!���J<&&�q1Y�:(��D�����m�+ۈ�~���l�䑲�k��IdYw��:��%�#�*,���}�y5h�~f�2��Ur$��>���ݔ� �n=�knЄ�]S��T���b��dSJ"Y�F'�J�J�Sʥ2.�.�Y9v���=�p֨�5���W��R)ĖT���scq���qRk148�5����QR<v�a��"��K�/O!cNJ��ۧ6Hs����v*�+ih�=������34�?{���!��[)�I����ic\s�À��"n�>
����pm��}b?����W���P�7�<7kab(�|V�A���#ň)�z�䘢5)�uO$��Ra��mK���T�1ʘfㄱRS�gh����W_ƞ=�x��?a�����YI���ڊ�#"�ŭ�&}��8r�^�57}���LC�����{�B�R�ŋ��g1>9�Msb҄`�B��F�AxI=#�������>�gd�eP�؎T쑑b(k_u��D?+�]dhZ|/��n��y��84f��T?2o7xr����G���m ���OE@���Ei��?��E"�m�kuZD4M�?4�uꙣeܘ���A��>����V!n"�j�iۥ~��i�mI�>΀P�"�E��m��OX<66��k�>)��Ҡ��`��	a�I����&੧>G�ī�%M	�ݏn����]&���9H�,1Y�t/�/������wE�Zc@)�����[��z^.C��CfL�������bZ2h�\]�*��,S�7:>�&�I.���'�~;��9�����W��h��/}9K��@�.G��0Gah�Q
�.ܨٿ?��S{R4s�1�H�~�1-���X.�y���H���Na�k;vD�M�.H�B$�(�s=ީ{��`l������˨^�I��O��zf�o"i�V�ؙ�At�lSr	soz�vTiϻy���"��m���2�1�H�_��HһLSUf`&u�(��0|?fB$��LQ�9�2ߜ�йSF^G�+$�&c�I�EG�0Bq<f�>H�ᗮU�PE�J�qz=����4�����x9�X+���vϕ�*q���nM��cWMKPV��=��)b���K)#��A��l��Nɴ	E�y��#������^*�p܈�`c�Q���&n2���,�m����&�a�	EK;d��-	�r�B�V|�$�P���>bI��v�{7�썚��0�wo��u�8!-4�6��G葚��ii�Cz�F���Mn���Ќ��4����3½���>�X���97��a�=G�o5m\[�D[w.b�f#��n��$�K�.F��01�f��L�ty]+���9]7P�/�_����H[��)kq�@/angzQ�Ǖc{��2�w�t��Qx�P��v׻-�� �Q��n.�Ʉ��ۭf��'���ϵ�/C������IjS"�8DBP�����X�ZPetm��:͍K�|%Q�2v�;2�Ĉ�"��ȏ{[efy4�)n�����0���]P�N�O������殧�{w�j��vk�G�/J��L��\��e	�3۹�0��*��7��ݐRU�F���A�ݦ${R�iy��B�ػ ���*
E��+�r��E���!�̾&X r	�o2�S��,ߤ��*�Kԣ�G`0��� �VI�mbv�N���cwp�߻�ӻ�e��c�;1k�}�hgmT���T�Y
i&��Vi��t7�Zp2[�N�&�Zm�<!3�n��1s����4Y��6��̵yj(eC](G`+�5Y�(K����y/� �k˿̴��˫��1��A��5g3L�k��I�)�z���i�z�I��%xj��c��v��y�/v��N���S�ѻ�)��K���R�/L��
JS�8���Q;���'C� �+:�
����&��[�n
,t�b���M|z҆�eP�7u��֪�%��%p6`$�|$D���fCn2��c��,-�����k򦋏�<|/SnA���p�0�����z?�j�`n�������T��/��_l4�i��X��3��{|b�X{��=���>�_������(���2��c�s�x�:�7�Q�\��卲� c!A�?5��o[W�1@��T���Z�:��<Qю,YnSC�d����٦��-�dJ��q�C�x�q�­��H��z��i��n)����K�8�Bm��-K������1݊�v(��.ޟ,�iZ�&B�La��a��f9{���-�N�MI��c�������/�\A��а,`��Ȕ�|�Ԅ]���Ԇ��:j�#���O�_�C
���*�*����P8�����e
��f�#k��U��2K
]B�Ծ���;]�0u��y�{��o/��@s���b��~��&/]9�V\�ع��ƥ���}:�VƸ��3�� �rr=� ���WH(������nGOc�G���K���	��(����wd���8M���M�q��%s*���Х�%�+�"�J���љ� ��⦄�I;� u�*O9�|�>�4��t��r��II�4.$�D�diV����%�=�+"���҃�mB�DN�O5#eJ<�`ۄ��/��f��� ���>YQ�L�l7Wt�ܠ$4���o���'QۚG��T� '����C��?�?p���d�s��,�yg_cY��ɴc��󛍧��m.�.�/vH����$~���x�3��"X^�~� t�d}�5� h٧s�V�8�G��u����i�L�o���e\�AR�H��!�&��X�6�[d~���4���{&>]�Z`��b�6������9�PaPI�H���DfG4C�$�v��O��E���$�+���ɟ�	������x2L���m/��o�a�c�����p���a�"��:��Ј��ztV�OZ"u��x���RG_\nk/̬�E�"Ad(sڥy-C�ܭbѸ� Y�&
b��ja��!��U%���/#^%H����H8���Y���ޒk
䧘b�1:oÈg㊍�&�x"�N��L�Ѥ�<��7[	`�Y�65Sސ k��h�Y��Q4#e������15u�{���BuYj������Fexő�V߄J,!K��qð3Cf�?1e]Y2L�i@"P����^��C�k��[{D�&'
(�h��<ޟ]�u���Ҟ��b$�`�Д�K]\�0 �s�P����t,J0-���5q�Q"���k.��H�/ė�0_\IF|�N�kh9��'�]�q��28���z
#���Q��pD�
���(T���P����~�[ߊ�\|����_�H���0J�(S����:ӇǏ��C��&MNS��1}ēO��8��,������[�u_^{#����<�U)���A;۲ui��V�h�K<���)Ҫ�V7�$�$�ڮ�/K�M��o��;&�S��k#�D%�����HmC����&UA#i�5�t�È�B�؆���0�U�8N1mj2{`
E��&mT��5q�R��˟��?��GO��vq�?�$��{�^A�30>jc�$�^o��+/��D0$ſ �r.Ob�b�R(A��l)�P�DH���BьN��8ddH����M�%В|G��̌���f0��d�$%�:�0Y?(	̄QJ��V�xU%L���(ٮ�b����A|H�,������	%��8m9H�(TG������+f�/���&s�eV��B�fM���quaAp�Ժb�\�W�W�>cw�Q,vr0�"ȾC;�Fc(@y��w��4n�B�k�#�Z��B�r��s0:�E_E�o�7n"�p����:u�����Fw���(N"��2a���hg�n"wv��^) }=�"��`/�]
9��e�c(�4$Q���X��tF�MS����UF�T��(���3fOgI� �4-b�(0J�_������R��m�bf`fPA������k{��uD[��p���^`z����uX}��Ml43(�`l|������І�dۨE69@�
I�ۅa��r(wְ�^����j[���"���ob%q��Ց�8�8W��4sy]��4�T#���Y��4ֈ%���Da�.;�viK�U�ʝJ�N�ҷ� �K�$�2�L'�/�W�1����hK�T��V�%i�+��8ǧ&��I7���w��gl����3��ъ�ȍᵫ�c�tN�Y<��������67y���l��Ҩ��m���?�`xܡ�*��a���Ը�� $$���;�@HV$�Enܽ0F%)Ft��o��wē�D�����,��}��/1�c{f�F<���I>)��$�����k��*@QrR⯬�;� �/�8�([\7O_Р�O^>��`��	��ї��E��
�!�x�q��/�/ɪ��YI{�K���B��~�>2B����{�]�R��K8��ƌ�����"I����t�K��ÿsYck��`��Y"�=+�-$N]�*������F�a�E���5c�)a"l���W%��$Aޓ���j�a�Ů(��qʢl)��8A���E��!L�s�����l����w/�>�ǞÇq��Y̝�5�W�v[��4���Z.�u����Ĕ�y8����[�x�ډ�:YFB����A�aG��k�eJ9|Y���F���9N{�[��VFpQZ�L��#/��+��{cЦ�T_��A^d�-���C$B}�8R5ݼ�gM}ݕ�8@2��a��7CVHk�q�;����.ǭf͐��|6+�;�_��y7�6=�K씝2=M+od`��-(����M���o���W�i�ju��=���+��ހK�����wH:Yitv��OcD��`�V��e[���U�j�1�U��ho�K��*�����M$3�� 0��-˱(�W�A7p���k[�V���0�)���?�޿x�&��Q�;��&>:R �?��ҹ���X_�a$()��ے-&ď�D���BaC͘ -qGA�v�;v?���9���Ԍ���47��c��U���F���j�P���П�x���S    IEND�B`�PK   T��Z�Bʟ�� Y� /   images/8b28e7b8-a93b-45a9-8e01-1e8c89928838.png 9@ƿ�PNG

   IHDR  y     ??�l   	pHYs  �  ��+  ��IDATx��ٯ%I�'�����v��2�*����k��K���� � �x@��'��zC�G�Z��Sk$4��̴jF3=�PU�M֖�[DFč{�.g����>3;Ǯ�9�fUk�C'�Y|177�}�o��������տ�����������W�w�"@u]R�T�%�3��!�<����-Q���k�G�(�K
�*[���A2��ϩ�%��싿�ùx�(��-�t|L���/��q��}���kt�<�9/�qpp�mm��榛L�EF��ʏ�u^�e��7�*�<߫�"������� �W��M]E�p�m������͠kګ��W�"
��j�Z����`TA����X%u~]���E���AI_n_n_n_n�/o����'OT�]����ڧ��C�8���ϯ)M#���������*�i�dZ�R���g�+~[S[�w���j!@�![�uÿ��i��o���|�ǉ�y��S�^ �������S-%р.�L9-��ʳURT5�J�pt���a�U��¡�뚅GP�^��_{޺�<����jZj�b]U���.���Ni��+�8(��Z�*_��z�xU��n�e�.�d^�O��|�"g����i��*T�/˺�n�����:+�L|j�kZ��E�����/�/�/�/�_q��������%aB�Ʉf��;�ٳ"?���2���4�fj?�T� �/�*��	���7�'>��CX@H �;���:>O����AP�� ��|��'}���E���7>F1�W|x~�Z�|���5�0�I���1���8�=�r�Kx!_��z  ��)%逊����5Ō�y��c����m5|M����k���J�ҜO�SS���z�$��`����Mu~�h�O�W�ᰈ�p�,/�G�&���7����"��l�Γ��_��I:.U\�Ir@O����_��ш����eY\-��/�E��o?�M�|�}�}���t������^���~@�#bˀ��f˜��ɬ'���7B�;�.k���>�~_tT�8kE7�"�\�P�ր�����}�S����%O��@��9��`> �|Y������x8 �����e�51�2�*m.�=�W��`��3Q��h:���Z�q#��9��cU7��u��G!�� ��`�M$�{M����DX��T�8�)j�nѝ=_4��^�a����٧��8=}����x]�e�"����y��_�CjW����GӃgFo/��y�?��8�Hͫb����|5~�W*�볋"�OFI��i�����i��}�}�}��+���i��Gi��/f�!MF)-o������� P�W�60�0��Lcl�-�cĔ��4�1��몡l�4�Ä�w�s���+  gl����<?��:�����ä�k�>pY��'��E]�&�r�QWw�������95E%f�NLE�����h�P���W԰&@�{�R�e�����=����.WT��u!����5#}M�D��#�������./����-�K�9�aHk>�Z����R���~vvF�N��l᭳�ø{��wʏ>�$X��X������4����,M+֬
���*[f���q�\ϗ���բl����88����O��5�����4��l����-O�ӎդ�[�_O�������R�t0�����ng��nz=�>X��o�F����{��^�/�Wx>���x�������������������>P��w��<&���E�O&C?IJ���o�מW���'e98??��8��t�������駟v�=��?N>��1�a�@3��:91����r��Gb�������iGh
 l*a�)�-�,P���@��VUA��1N�!�f� E0`y�A�p��4�E-`���ū��9���w5_��%d��0��,wk8���x1dq�,��qSR�x0�К5���6�1���8w�WP!��~(��σ�PT6��>�Z4!i3�}��L�А'��k��Ǧ�hY,h8���kiCȍ�L� &�ׯ^����b����L���t�5-ON��'îfA��Xs��<������3�Y���fU��Y��$�f����J}��M>
��n��󳧋��>+�^��VEޝ���R��zX��=��o��EV�ه������O�W�����[O����~����d׋Ey��i�_���Y��+�B��K�Q�\^7׋yy0<����o�_^^<_������qx��oc>z��������?�i�Ϭ�F>kV���Y�����7��:���j_�x����]^f�Ç��?e������owV�>���]syyY���4���w�#������܍�_����P44y�ϟ?gm+W��~�X,p.��k_{��>���f�� �=���5?�&ϝ��h��������0��;�������㏹�S������ٳ�'w����{��ks3���fg�lVv��#@��b2�a>�^�̻�����Jv��!�������?+|�1�&�E2��|>��|�j:L6ޠ����8�9�s�����˒� �$ڮ&���^�ۗ/�e׊��0��
yU�A���yܷ<����8o��w|n������O0_Ym�wAt��0�X��4%` ��|7���x��Yp��}�{��[��H�2��� �1Q������EQ�|?U������֫�u���<y�^_g��d~�h�G��;�|����+|��=�>�V�����|���(J��
c�뭯���I�:�drp%y�dYz�~�쭝_/����?�~wzx��.���]�4C�7�����A����Y���g@]�9�̐���`D�Y&�G�y���q��|�
�����5����`:����͙у���r8�2 ����5^-��Y�$V��C;�9���Ӷ�4��@yY,G>  q,�7�� �(U�2���Q9f���1P��8Y;�B��@��}�}&��V9�%�m(GE�A�i �}0�UW�����	چ�L4��UV�n�ܶ\4�0�����Z��3M%_s���|6g��1�DP��� ��@@�}��k���7�-���яQH H��8:��x8�B��#���㚵�nq���GM5Hx��]ÿ��AS�][�����	��kX�(/� 햳������0��$�j�u���z��IΓ�'t�@���va2�)]������?�C�<����D��]��ɻ&f<5�F�9O�%�����n8������(\��e�cd��~p0���_�R�7�����W<�ʜ��ѣǗ|^��'�'��bzxxrpvv1n���l��LƁ���0�NӶ(�c~���EAP�y^D�<��u^]�%�w�Z�y��|�,f�&�B���r����7��b�)��|;�����f b�r��o�˗/A�0p����'.�y��ܙ|aW7��[om|7�'ꢶ�f�h<R�:F�a�ʋ2���c�x������ap�\M���{�x�u���Aǘ�v��]<4j�� ��#1@������L���^[����N$~U�~��M�Z�A�t�V�s��	���B�*�EF����?�<VA��ge=���6e����m�����,��q�D*�v�v󶠭�bP-ː�Pכ���B1Fe�U�q������`�Y����gv��Z��n2�,|�x0���Ϫ�t���'-����Ȳ�7����y2�����<��c훟Sv>�m�b�o�i�y~�Ayxt��q<��v��%m�6H	��A豰Pw�������>����~���gr>=yp��2�S�8���A4fp���D�W���D��L�-o�����^13]-V��rh��>`� {0{	�d�/��w0�N�$c����4�� �����tǰKyb���Fi��p@O=`�e^�x���󈁵��a���1���T1�G"XQ�S��O%KݔL�"]����J����b�4�y�´�s�&����C�!<T�A��A��Bh�5�Sa���+b\��j!��X��ba
k��A�����5IX���G���v�?T�t�`}u����J��"�sjYz3ns;�rS5���x>R���B1�*���
GT�X��4/�r~:Q�V�+0�����,x�i1�Z�6QSr�th-߿�X-��1kK�nt����\<gaz|�w޿eA�hmO�sp`�i:��B7������ۃ��σ��@�C��F��qQ�!�/��1ǁ���- ��D�Aڲj�6�Fa֠m �w�����7$0T"�m�De_f�i�����2����3�5�֤�29� ��b�`�v|�0��5u�Ʃ���C�_�������xޗ� UB�c��,&�D��V���t æa��y�I�ǒ�c�dݡ=|����*�s½��p��<X-m�[g���#��ca����3�g���29�f���@�7�y0L-�'*&q$�-�yß�}��w�ZO�}H�"���>��P�l����E�����?�~;��0���yh������hV����	�e�˥7�NA`un�^��S�ү�Ҍw��[7k��}�y@��D�3��
��JGv�4�Ě��@_~G�^�w����~�&���M���V���೜�}a�5����(�G4�b�yT�p�&��ϗ'�Z '�0S��y}�k��*c��`����x�� )ybh���+>����ӵњKe���,��,xx�z�䁢#v`��% ;b��	�� �m?�0p���&����ί��"1o�5�>A�!��-arR���	p��R���8�k6Ҷ����lu� N0���W�y@�!$�2��������ڜ�d+B��|f�S��b�E�S]�t��D�g=�S���F-0ER�=G
�c�a�C�=�.�S�3�m��^����L�����̮(Mqb�OTJF�<K��b9�� ��M�Ȃ4��fP��a�秃�}�x:=D���B$
�7��x0�Z���������&�!�\���=�NO=F0�[&	ﵙP��c"�x"�,$�@Q�`�6���u0옸ɹD���<��ad��A�M(q=Kn h���8�v�}ƂvŚ���0�±��k�C1_2�˜�uX�h�L�ye��2G$H�ӑcE�������.6��l���KX��	c��p6ܟC
\����SD������|��ԉ��0D�Ú���l�X�+�Y�g:���=X3.�
��m��g<�y'"�Jn�Λ10���WpS�/�o�_̡HůȟC�_��?n+ڤ�i��Q|��_��F��bc���E�{�cD��rӷ�C������x����hk���;A������W��q���?#4f���!DȌF�fE�����Y.����97V;.����<�f�?�9X�<��$�Yf����dE#�/�S���Q��������L6�],s�a� *���,x �'�m��A���!?LL�kD�\�:��dJǇST	����zƃ��v�DHF���Y2�A@���0o�MH�����k@_.3X0�͖b�a�OQ�pP�XV&TƩ�7����I�m4��g���yR@聲��(7����y�#AJ�E8?�V��h6M����Ɇ�*}N_���6������_�Y��DRumD����G,�;���A,&8�/`u�j�g'5��q��������@���c�@ U@����4.xbmr,��/��8�y[��p�f�
Lӷ`�}q~����c}����-0�`��-Ix�V������a�#1*����FxTU-@f�޿=��V�6��w����M�V�v����R�-Z_��!�vm_X�`A�=���y[��m�}L�� ��C<;{-VC(3���g��+A�9N����!�<7�<p/���m�ٶ�޳m�K옶�V����}V�v��$�n3l[�=c2@wly�BE�����<n�ѻ4Lr�<���Ɠ�����UM�EɀI���;9�0�٦I���(�J@*f���&)����Ε� $=k��H��̳��J�@ZӍ��V���� O:L6���R0�F,>d�X|�#��f:X���trx@�;Ox�s����m�p!��R�97��0P���-3D��  %߼�U��E��x[�f$� �\�y��0��'f������{k�Z~���X��0�I��Z�ݴ�&�C���8.�VM���"YH1�����y<QY�f���Al&w	��2@�s�[% �8�*�	k�$��ς"��|M�n'�|��~	;!Z�ޜǲ&lvl���	Mݚ\�D��`�u;`B��?���[��u|o"�H��̄��>(�ߛM�@�9���0܆�J[Z���y �r��з������l7y�]g�^HƎ�l�sY�`�� {}W�Y���|ۧS�>W+�����N�~1?Z�+�6�o��p3�g����>"���� �+h����;�z���}�YmD��ˋl��ʌ��=ڗՈ4vn�Jk�o��8W`��-�+&&��P���?�<Q_=�t8��_R���G������b��{8Y]Y h���Pag�k�@��O�Wg��!�+�~xu~-Sذ)k�H�Tc�ά����F��1a��~`�i�0(�)�:��S�*�Y�0��d��ɲ�d�P]�4����H��>���j]K���!a��v�I)k@��<�-1���	��t��T�m1�0�Ϊ�ִP���t�$N@��Cug����� ��a����%Ŀn���e���~���va���s+Q<8���`RW�Z¼X{���	�̢kC���)e�H_j�Qd�YP�Lc�e���y�9*�������`a�;�ܿ��X��[���O��U��	A�FU׾�x��T;I�g������]����@�7�d�+!|�=�/{nݔ��n.�t�w���<��fٹ\� �v�yFK7f��z���V�؎���� ���k�7��`�X�+��J��k:�][�g'��pK[�[�vێZ����[��}�8ƈ5O��i5{�����{6�/�pow�|0��y'~�� QW��W���tH�!��D��^<�ׯgT�T�+��ɐ�U�߿�y[aH˕f�����cVUF<)-DÐ�IE�6 �1'�pCp�)m6 ���Nr��L�ذJFcL8��
�6��0��fU^��/P��҃	�o�׿ZѧŇt|zB��)���
=���D�!d��d�t�06l�0� �����"
�K�jEu���Z�Ё6����d43�Y��4M�鉙i�^k@[Q����nC��v�X5WzC�o�xf�8�
�о�N?��hNx(�L��ّ1��F#����&�h���u��1����x@�``WHF(�du8��&�*�����L^~n�5&o� ��~��Lj�3�ZV�u�9lL��0L;��YM�2�U.�2m6$mcv�c��2��U�u��fg.s��HXF���g�9���Ʀ���MB�C��@t�-aR���`�m�#�l{�o�'��'�zx�?�X�Z�k����Z4-��.H�>�������ע�'[?�j#�@.�g����6c��w Mh���x���
i_']B�����g�M{o���������y��)���5k�v�bxXR����ִ����e�tW{+:{������|�ے����#f�%�����Ӄӷ����矟��a�)��y&��Fc��|���EB~��t�, v��; �!UG>��Bh���b���-��`�|�a�H&����?���h%&�+�R�/B=�o	S�b㩫���y�Ň,�Z��-./H5�8���'tu=�E��}�bb���Q�V��M��R4���t8%��4�?p�k��\a�A�Gp@��X����ھ/�2��Wl[k�4c��*1�X;v �t0Lha�i��pz��Δ���6��NB9?�@�NL�G��ؘ����!=x�U��'�(#�^�F�0�3�?�ހ� �0�2�wm�C4�H��;q���,� o&�kيz���:�t{�.�[#�.�vY����:����.�{�d�
���5���9�� ��^Y������������ƴ�����n�m����7���d�^��Z�c�a��g���0yW���-H�M��o�B�e���}�j�%�n� O�?�5��p��IB�yF[s���cǁ�Ķ��m���f��:�]��y��[�	B��
Xh"'''w��Ƀ�`��:����LL[�X� 8�����LT���	�;���b��˗���������%�>��޻Z���3���Il�h��u!�|2PRu������P߬�, !��Ǧ���EBo���D�r�G?�J��|���fDb��������ǯ�@��J�'Hr*s�F"v)�k�Z�r�x��J:���M�$ ���T�K��a�0���C�!/�T�4 ��J����H�l���$�v��& � �ƾĹՆ6҉�M¬��<��5�Y%HB�5}:m���B��0b�U���h3JWo�x��`U,P^����#�o.1*�h�0���4}�M�����)�58�`m;Ķ�B�Hh#0Y�@b��f��-�Ԁ�3�=o;��#�Nkco��]��85����m痝d�W���NTk�q̪��\�j�c�t�{>}6�j��bí�Pm�koݗ�;{?nԋ{��D״�&H�]P�3��-0�k����Ld��.s����c�6���c�l50T��k�����c�����@��SƬI��qhB��L��X�����~�o�ٸ}o?�mk�?w_wk*��X���L ǝ �駟tq5���`�X�"+$2�����w,U�O�?�����sz��o�;�G�*�������6��g��G�4_\� Q��'�*pM �s�6A�+� ��l���ׁKB����.M&���T�z�LmlMJ��iۉ-N� �u$I� ��)V&�#���ZA2ވ�qzѻ�i�X��Ղf��d�U�r������x�w�j���q|2���c:8�p�uf�@�`�0OA�[�0k�!����z=�#7������׶eBo�X���V+A����iFo&�9��A#]b!ߵ�W�k�A'��\R{�=�sGSz#�X��:k���Ln�� }c�
X��~�0&�=�
	g�^����~%���-͇�ܱ*wo.�f2 |P�9E�NO��2��"I��N3����[?'�،ߡ5�=�=>��	�򶟥T���=AP�7��Ξ��m����i��s�M�@'E�5x������m���;怣��-����3�������fs�c����~�
�����i0|�M�u�lϩ�3�� ��h�h=}�B�x�dMS�P�$�FQY�w�Pױj:47�7��%@6���E뀟2�3~!�.���tǶ\ܴ��{x:��łv-��
�؟�xF��O����-�����Q���S�?`���{�oS�l�XW��/>���A�<9���$��gg�W��|��I;0�Bac'�%�P:���	��o��o��o�-�$�ǴZ���?��4�e�T�1�O���T��<�bҖ!�^�2�e13�a���X��PL1y�qrz��G3:>�4��+n��Mt�COO'��{t0�s�m�&��ԣé.����
٨%T�W�<����D�{�C��R`+I�V��VX�0v�cxa�w��,p����i��c�A�Jԣ0�Z �=�m,+G�*�Y�d�X���#>%hz��'�!{��VEʿ�4�5����:���e\0#h��M֓��t;l��F��*��c��x���*ͮ��i�vsk*q'����Q��=H�R-�1�|�<�³���	�8X�8�{Ѹ*��q�:
`"y泒�'o�W�9��ł��`�3ciyC��6�Z�_Dq�)q��� ��|w�=��A>P����܍��e�qLV�������u����P��>��m������G�|v6���P�d��e��5�<���`Y�,�Ll߸���HR�Ѻ �_�j�c��[����hȧ鶑< 8Ɔ��ي����Z�WL�3	���}���q~��_D�@����5�+�P`������o�ǟ|$���/��'tq��7<�����Ϙ����'���������-�����h��x6_���33�T��ãz$�;}kDO�:��$���t3������ӧ��̖ci7J`�!a�`�2��y���O
!�<�S%���	YQ�L�{��M%L*eA 6{�������^B	��G�M-���T&�/FuC��Đ�m��W�~��t~~�3{y�TR,�gcZ�����ہ�$�L�Rw�v-`�B1��A	0��/�,Qޔ�,�nk�$�� 
�V��JW�d��zQP��aؽ=��g�$�UL��bM���uu�}Rѐ_]��~y�ט���ph�n���(������A(B��T�7����z���w3�����cm�2q�6���*�c]S� [��چ���˪��"Uv���&�۵3[ߚ}��8���m����ms�������}㆓��v�Q\A㶿o�p����Bض��7�{�}Aa�"МOO�7m����o�е��0i"Um����y���fF0r�k�k�m�;�Z!������B@ �����D�>�ec+��\�9��Fwl�������_|��h�fe����a�`G�����g�h4=`0T|b�7��ӗ�/���(5}�[���׾�\����>��a����7����}�7�'ԥuqEW�7tu5c�^�����C�v*$']S3D ނ~�����9e+m͐j��"���ҭ�h4$V�H��3Nء8�;I�AV�h5-�l�!��#��P ��rf��� Y3�S�D���Sue�����.��ĕ<8D-�����F��c>��`� ʬ3Nt؞T��̓
��3���D����6�Y���a�A��xe��6�(��$�-���f/D��&t�0 wd9|q���ѱ�2N����;�~����_!���2y[�[*�$����싩C"}H�je2z�I蓍��u����G'h�Z���N�8o"/���u]����
�[;G�pm��?`���ݪ�v\���tnk����
�]L^���na�s?t���m���}���:���rA�e�n;�}n;B�L�h��Z�]:�+|g��Z�An��.�h�/��wY_���G?��F��\:���\ߚs�c﷉}|l�e��W�["����[d4pE�����6�����܈&x'������<X���7���(�J��Lt)F�7�` ����z��_���C�+f���U�:iQ���G'�a"�����矽���K���QE�����{_y�����t6$��C>��)[^2�������ё�B��X��l���A��	}rГǇ���8��Z�}���P Y�!�a�ܙp����t��E�>�׬�53��)p���\�Z�g//��ԕȫ\:y��,Al�erm���6N ���IM�$	D�"�(Q�٪��ԧAYc�e���1V���\�Ͱ�V `����'J�d@���x��UM^�sġ˂r���!�48ä]SO>�F2���`B9�D��kJ2��ꀖŚA�@8a�6N�SCc �p������t�q�"�QA��MT(��r�ÑDz�F#��-��$�~��Q�,S���&��y�F/�ځ��~炇+d,w����u{n�	�Q�;���F�g��w;������2�}l�J�_��D,��[[���~\Vl�w��{]���Xs�}&�:W�F[����7�H6��\�j<V���׭9�2{ԌA 	����o�����8�fO��Y'>څ�!�$����Ƃ�$F"�1�Nn9�W|�+&ٸ�~��M�6��/���������N���N}��߹�n>U�!ps����10N�X�<�[f�W�|'|�}D���O?��W/.��z�=<�'��@�>���x����&í�������I�R��a�i��t�t���c�nѣ�	?���X[!��lLO�0����*V����T��T%&8�#�cj�
�<K'�r`� �;�/ϥ�q4��0;�}z~vM��r��i$l�h�ğ�N���)�<OY8Fr_`�g/_���nh����R�`�\����Xz����uHI��1[���Ui�-,�&/��Vg�t5Ѐ5�2׌k�$C}���m�)4�Q(eVނ9��MĐҎA�%b�K]#�8�y0�M׫�|� ? ,�(&&����0�>kN�h�(Ǭ����E]pO �D,���`��yЪ��ߨ�:N۵�:+رU�
�.�����-;r��kJp��}V�/Jb�LM��0�i�K�g�6��=���M�����]A���l�j�nm�>����]���#э�q�o#d��b�@���-���\ML$s��6���[MضŌ�J������t �P���� n��y+xE�4&��5�����!cֻt8=،/Tԕ�Ä��8M#��\lk��^�3-�-�8~=�go��vv'ȯ�u���/�������xd�0kZ�K,r!�q�@�b�MxBw�$=��G7�5:Z��jIϟ��b>���^���]�]]]I|�K������¼ x���ߦ�����1������y��{�P����TL�x��T���$jGЋ����6�.O��%Fq�`�E�֬���n����v��P�3�W�p�z�/

ECf�(�	�1b"Y
U�����\lۯ�
~�deF�Y�`�����IFc� w�1�ŕ��X����xv�
�FY�	�Fl�(��lQ��5�r_M�L��8�����^\IV��ǧtz|B�|�]�2��+`*�`��֮Q!vN���)�^~|������g�πOd�V�e����&{�H
8YU`l憥��\���.Ƞ�n�y��'h�`�)��4���F��D�,��@���.���q�ov迷�G\�rA�=�{�U7t�o��3�}�%�8m��a�oٻ,���
����?�	���ݬ��ߏ���v^s��嘰�D*�mS�:�����:�m�n�dVcԶw�n����-Y���f�J��8f�_&L���S�q�J 
���J��x�(�}ܵ�O�8zZ��� �ٳ�������^����?�g?{v{*fU�+��4����5���:c̀�X͸A�$'!�3��D {�d��h�D��Rb;�^�b��1���w�Tͅ����1#-+�E�yO��p�\�����0�<�0a5�ƆɆ!
�l��X��r�,|-��5`���J�Wc�׷ΔZ ,>_iSP�x�����%�.s1��}��x0`�p� ��ٲ�h]�2�J�=�Ӊ�!p�<�qU���'/�<��;�w�M0f���=�2::�&�D4.�K�$la�t	�#iL�j�Θv��A���G��+�Ӈ�$T�v�lTz��x��D���Y�XhR8�i����(���~,��#�-�I,QIX=�#sQ��+}�l@^ ����Zc�҈%��K��F�-Km��D��lNl�Ax��Y�>�>��b�n��&��ښ�}�ɺf#7w`�����=v�ZG�5���V�d?[��f����k�>�f�w����}˦�LZ��<�� s���ʡo�R�N֭�q��k�v��`s���]+=�� �6���k���|pg�����V�����zS�B�]��e(��s��@8c��O���3��!���_�����������^���F�ӣI◍�*I��!J��y��A� �1|��xn�Y�IJ�]IA���vDG�Tꥇ�ՒbEJʔ����\��}���bj��7�t�[f�c
>0�X����lI����/��fļ�침���������R�U$�)	�W���ťÈj�H<��3�0_�Z�":b�<�˫\"$̩Q��2H�Tl� ��Y���9B"3$��Pw�,٨�Q�j�&�/�V��L���$A!!J�1la/�f-B�w�i�tf֐P-s��ġAK��d�Y�X�8}�X�aӮ����|E� ҙr`R���WXm�m�J�@��+<h|O~8���'|-ؕ���`�� ��G|EV�1YL^� ����$�<:X&��e�!�j���~��%I�\��4�&(	{�,W �ق�.s����2#X�p�h����[�Ֆ��m�Yf���^�5�� ����J\sK�v�/.f�-��7׸[_�� �-b����rߎ��G�~7����9�1��.��
w�vz�n��־9::�k#m,��XXE��E�����[��5�X'�Dڀ�2�C@\^^�__�|�Z������~��W�۱�^���<
۪:Um��ٴeS`�tA&Ė�ysaV���HX��l� ��f\�ĎS��b 7ԹQ�8W�׾N�G���%��k�*iִx}ɪ7�[�c#vU�k�2���	������������G�������;�\[�6�|��m`��ŷ�P�&	d��5ڐ�NW�C��ǂe�f�f6�37��Y��$�d=ط�} vc�� B��W����Y �D� p�΅�G؉��1�K*���=!t�-ua2YʐAq��"�r[m�s����	��P���̆Q�W����&BņAJ:6x�#��8�g�5sKn�Y>���f�d��1�s��� �G$Q�8+���8��oY�	�s&2
TY���������W��'�K8��m��MW��H�7�s��p��d�f
wk��e�����m�뷫���蛝���}����b��
2�O�]��������3�[��Qh�@��~�sب%�T�M��m�����
�l��P۰˕X�ͳ�E|!�w��g����y��?�������Үm/��7��L��i�xIОs�nLa/�|��Z&J�.�+qޡ��p�PŠP����<�O����Nk�����zL�}�=��B�޿Bb!C����ӗ4���D�1�M�E���lE�k�`��V;%��<��<Y��[��0>M��4i�F��Qs$$�/�>#�H{µ�2M�2�Qr�E��bsg���t�����:O�"1[$�:�Y!4��V��)� ��t���܀�T�$�����UJC(�l�n��D���<��mS�������{ǂpڈFd"z_m�^��Z-*��i��&�HX.�&��rA�7�zz��1��v���.Ҧ#P�YX��e�$��)p�l�y�D�V@�kF��ٺ ��W�N�i���{7N�����پ����׶���
��9ݭ�m�uN����ic�u}���>����<��������.��5Q�}v��.mJ�v��6�҂��jMVk��m�^w�ۮ���}l�nB��p����NZl��D�C���!+�z���Ă ���5O�x��%ݱ����84j0��Ԝ��&�|����W$�>�̝$�s�����i1��y��4��FnfE�^��1M"��U~����/$N�f0[��dK�nۜ��i(�#���Z��R�`�3�ep�!��ֵ���^^jS@WI��7��<PJ��_�]HѮ0�(a�/�J�@L1d�d�D�\�f��tt|�K&c�� ����}^'#],�� $���%�W���m����䉮6�&����[�$QEm�#O�b-��_�����P&��Ȅ�`�ZS`KL &i�7u�%����D�uH�IDՐ7f��I������6�x,L�u}g��G,Llx~����)�+�lAކ`n�/����f�V��5�-��͵[`�����n�ᶗ�:�v7�LႥ��}���}�������lkؿ��Ǯ{p�kM;�~w��l�v����i�6�}��n:��v�bWp�}*���ܥ	�����[����S�Ygrx������l�1��W2���������g��?��?Z��^���F%]�t��D�O��� n[�J��`[`�HDf�؅���_�ʑ3,
��@�]� '@ؿ�:���'�>�E'����9]\�iveja�1.���y3�W�`L�IB�Pы��M-�NB�FT�9�p%K�n��Ţ�,0rx8�l��	%�P��`*BbV�x�/��"|Lu�������S)P�cf����|U�P��马w�e� r#t�W൲�,��!zf)��Q'�+� �&�M�b�oc&=[d��u��g/:	&��,E���#� �2�$�ҵ�rZ��G �B���{$��e+I�׉R�/  f�i؍����-ʢ����U�0�D�J� 0PF����ܘ�|��*~6�ۖ��(�IJ�xj-��d�����#�n��;�]�s'�.��5-���"��ٯ�������ݶߵ����{t��>�o_�����f����߱�ǳ{�/a��B�1�h�4�����6�w|���&��/L4 xD�'��3 ȑg��;�	f�� �W�`���E�K�g��Gq�^�>�)c~Jp�Aڀ}�ƻ�`����ܒ��b��c8�Po]�@����RZ�.IZS�����?{�����GOӫ�K	+\�9h���7��&K�-JT���<���Jغ��Q:x��E�:mi���.ڜ���C��ͬ��D�L�LY��F|�?8la*87�X��n̑���������_o���	�ćq.�,ֶ�d��t6n��`w�r�RPbA���)) jۓ���)c������<[�r[k]�S&�]�5 #n�"4���$"=ȌP��i�	B��6�#��`F�z�O5l���$��ȄB�d+˪Y �/O�U�ZS�lkjBf���'��r�����S��K����f;io��L�I����>0�e#� �&��@aA��L��mT��+xv1ž`���} �ֺ�eA^�dsk�����t�}}sS�}�7��q��9-H�%,�����#u�L2�p�4q_kp}��y�Տ'�a��ԚѢn��|&�@$˥&9�b$�����5�������6��?����گ�S�����|�#w��C&���,���kY���"�.3篽��vٌ���P�C���F|�9�T[a❩�@�� 3�.Ġ,��F�F�<���1k�Mm<ҍ�?B�ؤ�#�����J��t3�v��k)��grp��`u
AÖ��/Y��M�0 u�p� ��%�,`���_#Ωdֿ,���偬<�x���Sͬ��I��	e5����.VИ�_��p�DD�����q#�l�El�Q��
 !"�d�����=�?�p�.�T۔��2^g�lX Fj�L���f@��D-ab< kd�/%}��K9���-���I
��EUic�m9���[Q��n�s��lF���t���b�}ж߹�A0��Hln��.���&��]a���lWw�e�q��Y���w]�o���]��g��:�>�Ov�������׳�'���s,�s\o�s����o_���R zk���F���j���z[N9,���Y}��Gk�g��Q�xeQ�Ecd��d�`p,@��Z�	��S�*
+a�y�����WKYc1�e�9��!hɀ��YU����K#)l� X�)Ӌ)[�*"3�!
j18#*�s����\@��p��t�}�k�KHv�]h��J?r$�(;L������t}s���%�-�P/[���#eD0�5��,{-q�ø֦� ��-�X��6g��Ţ���$�ş��O!�5��M�$�6y��8��`S__�.b[V�7�v ���t��6�e1�F�B+��s�Ί9:�E�����Okj����ƣ�?S�s�ht�U��ם���4v]Y������Ujɗdkɸ ���T�(5�*�ڣ֞�F��Й7��[ !q��Hͮ��w_w�:[&�fws��.��B��^WH� �&#��}�wY�>����c۱��q��1��]k��} �����Ѻ9� ����42�������� 7������n%|��� �"ys֔k@Yo�����L������D';
2��������(��	?� N��C�����Ճ0Y%-��4����_V�l1�)���Wbw��J���x��#�
�t;::���$K�ӣ1uW���8M�F���J$\'I��m�2��|O�u����G��<ôt��U��|���Ig�X2�򋵇t���9e<�$�,^�+3���5N��1q��*H�դZ��$�>�k��
}�ZYʰ����ĳ��[�Z�(%챦�I�c�j�_�j1��dL10e`�D��e`p{
��P�M�5�+�$jͺ7�Si!�'�J�*�(}i'��y}��Eh �w8���_�{����h�?`�q�	�����JT��Dra��-i��J���a����h&�m���,h�����Y��!w�>p�����J��G��P�MP�T��b��b�D��ѭk� ѻ4�[`��oܾ�e����`�����ڧ��p����O�k���]!��o�{����9}��:P�$*����>/Y�NX,0� ��#]�c�q�.��U3l�e8�l{A�Ƀ�8����ٽ.2
�%����	]���#Z �HL��1�3S�P��B<�N�/�P_��U ���u��g�ވv��F|���^5��,��"3(X��鈲E%�1>:=�@�b�OF2����">�=��#�z��j�`	�H{Se���g4�N(E�r���� H9>��� �hv=gMFg�2̲�E���m���9?t�<���v4��C�X:����Z�� ,1f �o@�0<Ț�'٩��"���
� mV�9�����"jSl���C��8٤�oU��z��)�������ִ	NhD�H樬iH~ lbf5?U!�눢����#�VQޥ�,�[S��$9�dS�c[�!f�Q�����ͱЋ�~��-�9����;Y�����;iw%��G�_d��w�Ѷ�&�Y&߿�.���|���c�o���?�g�g{�>Cw۷���܂f?�?�Bbۏ�f�<��"q�y��͸9n�B~��6��>?$E���]�R�0w�*i�&ݾ�-��w���O��|�����u���Ϟ�����a��E��DY"��~+�D ����td�3�嘨�D5`�!��0l�DZ������RS�`����ؘ�qPG}c��iL��TJ���3	5
Bd�$�*}��8E���-7��QL���<y��}Xxb���A|D�JM����x���ɘ�a��Z,oh��>>S��"�Ӓ��-�a\t����@/x�?mYP��4�!;��2[wԈo��±Z�9��Y^�,��M�`�x2ބJ�!KV
�n��TxSmC��Bm��S�z��J;�!��Q��)M
���(�pI-U	��P�1�!����X����tNm�&�����m������WMߵ��ٛ���8��6{�}�ٍ�p���o������Ql�ۜ�d׷����>!y�w�cw��6�b��=�ӄ\A�?V_�q{=��I�M�rC"���63�n����d�X���|�C&����&`i���Y{���X�=�^�/�"��N���*�V� ݊�IK�Y.1�p����%���XQF���Za�u����#�LQ�U���UV��W4���o?�����RN+�#%旦YP$q�	�_�5��Z�1�� �lV�^$�q�����ĩ�5���Ɓd��|��xI�yC���_{,�F���s�b�k�J�5�u-���U�<�a���F$��m)�ܠ>:���k�+Y~�m"�����K�S�Y.L�yF;L=�ӂ�R�Q@H��,��l\��6��L�aö*E&n�ӎ\Z�������P�o�UI	���i��x{�4P��b��$��;ё4��1Y��	��>@�����vB��nG��2S�"�w�����	/�2o�ԯq�˄�E {��w�����{��eW�ڿ�ڷ�_TӸk?l�8@�̃�,������]�걹q�6ʭMe�&q y.���F��fo9��	Qm׭���l{A~89����N�@W�,��:�[3��Qd��vP�j��9T�U۫���<ٽړ�r�gZ��雨�Ҕ��$���Oi4dJf���S��l����-���t��aHcEe��赘4`�E���D��µ�5�"L~�������� �=77�t���򥯝�k��Kq�B阠�Q> 5|%����<�^uI��:�χ�ė:�>�#J�^�ՙ���e��Rr�F/����Uꨓ�v��A��,���/�0a�500�5�6ʤ�57uƩ,?h׈5�靅I��#�40G�'�U�v��?�1�R9��F��$�5� _H'K�Y�kKlf��-���1�]&�]6d�u_����ܭ�݀翱�/�� ���ns���.��f�vk�X~���?O_����{����]�9�>�о����>�������n����g�nm[��e��u�\�Y��W՛��nMk�����%��)w}���^��P���(A:���%O�T�3vLI!M���Ib� pG�qX�uA�Ih���뉴f�i( C�..lPi���)�茙�^@z��`$'c� �����5��C�Q:l��#E�� �Z���5q��8�Є]_/���qXh�$�2��$����3�L"J���ť�{C�`�����
vp��Z�$J9,�Pb�vw!��g�d�N�8�v5%0wD n�s�,�sl�(K0Ь[B+��	.�g%��K �,2��e0�<d�@����7�\���l Y�=X�'N����:�Q���9_Wl���7U(;q�n��a��zQ|�o�Kv���ؘ�}� �n۷�����3Q��vgZ~�m�9��~����>�� �8��s�p���p�۫�s�yN{�����q�Ӽi���e��m�}�+�ʾ�/�hq����e*��5�X�w}d���vX�:ﺬDV����|2H�0L�U3�V�ˢ�弡$h�T3��4����Z�&U�������lܰN���LE���۲*��{c՚�jNY>c���"�X)�Pb�kH6�@A���a��q��^��k��5��j�k ���V���Ka�)ق|=����3�=v%+ɺ�bׇm�A�K��e
aԢX�Y�@ �r�";���Y3d���J�L#|R���!+E���	��ņHnjSF�v�J�I�� ��P��l��Bh�ĲZ���j�����k	?l�����@-�gP�'`�� �%Q+�/���+m���V�P�h��L�A���g~����,�}�����;~�]��N�g��}�1����޶�8��|v]�p��w�.�k��k{���1����N���]�֯RjAݖöa�ve+��m޴s�e�.q���(|-ԫ�o��˲U����W7�|�{�UΚ�8�#]v$��<�eK�� �NSA��;UI�0o�sHN��g`�漭
Ϛ�Y�0�¬+�P���7k���T�}�h:)�@�N�BYpD����m��Q�� ��Ĳbq���vn�kD��Ğ'�CC[�X눢�X�\K����65J�vk�4rx�����.,&/<xO�zA&|�q��$�U�<c�	e�#�ڼ�<_��t���%zr/���&٤)�T@�E����Ap�6fE���i��LR����[Ԗ�H�B��BB[$�@k6����㉖����9� �Ǥ��>��Ͼ�/���,v�-x��{?�}��{~��;����\��:���i`�y���_̜�=����}��2�.癵vk�ۺ�$�n����9�y��׮o��q��`��4�-7l��Vx�oE������>�9.?|�����<[�� Q0�{+�UyMQP�b���Q$�)�5�4xǔ\���7VP�������D@2���t|0���Q���RZ��G��P1�8�#�� X,`�њB�n�'i�j���DI�z-���$��R�f�)�춬�j���;�ڱf�y��	�j���SHR��=�׶_5:$̗gL�J0x8�!�R�
|���< X �p �fc�[z���H�t�VM��[26{G���L��dh�>�n;�z��W4�� �|��o���ᬟag�c5���[<��ӦS� ڂ�KJ�uZm߷�S�ɥ5��q'۾��M����n��9�����+$���K�M4v�]��뻾����m�wk�x�T��m���1��Nѿ���݃խ}����֮��g����>"ᮌ��f��6����i��&o��o���D8D�X?�l>����|��o�<�� �z~����ɣ�c�YP>_1��kZ�[J�V���������*o� �R��>��F�$�J�2�G�[1�p�h<�yTxYJ�R����a#*�y(��L�\�9��c~�F�6�t4�s�d]�Ry\:5���IH�R�I)a�-fk<͊����[)i	�b  �Jj]��k����+�/�4�ƀ���\,oWK�z��p�`��O�(�P"�pAh<^J��F��0������ �jYv�٘q_4�!� �}��z�����[-lHiV���Z����'��!	`�F����&�{�^E�hyr�<|.d
�ɵ�͹Ȥ*i߯I�Qo2�}��/f#����$�I�����A�������ڱ�ix�}���o�߮��{���o�m������'�~������m��i�߭���ywiz��7j�
jӌ�R�c2�B?��#sNI��Fb�.�.�/����;�O�m'��q������<V圲�k�ϖ�e�8,�(u���9J��;̍M tX�Tl͵$!T�J/
�P��x,���7�,�ET) ?�U�s�S��	��@|��D�����e5*|��׺���r��q��Cb�s�����+ߕhZ��SX��D��q높����K�Q��b��y��}X`������E�I�7�L�$R�`w����S��d�B�jK9�%�2y#��D\	á�kw�p�Ĥ����8Q!�$3TL7���5����@ԙ�������Y�Cn�IO�l��<��o��C�5&^>ҹ�b�O�!�#] ͘l��ئș�x6�t��~q�k�L��[_`�:�q �2�������������*�����E��.'�>��/ێ]��om�v_�L���&o�u��XS,
��e1��q�Wy�-��xpx0���g�bE)�z�l-
b�sPӑ���;%vit�+��D�v�{(�?��xy�NM�1�`��ZT�8��-�ĊQ:�N(�"$6D�`)�ά�,+&��*����"S��n��L����y�]@��\B�D8T�>`TDdKł��%��2�F�T�[�lhu�r���Iq����;1��YX��[���t��@������HydmZ�c��q��\v&~�ļo��NB4u�`cq��V�����������Й(�V@�ձ�0#�U+y���p�$_ڎ�8ȈU�{�F�:�F�R=#��6�_��U��>�`����D�o�'(����>�w���<�luKN�+m���� �0��H���C�G+ �sί+��������I f�	�'�O��׍.^=�>���0���\�V��h2���{��P� �,W�®>` �OR�Ʌ��YƀX0HΨb@��	ߨ/����,����T��S�cDi]݂�b�� �_[�F#�T�-�m����BeQ	�E���$.O;� d =�̀��y� ��� ���KQ�DKht��pľ���`]��l�/�.��O���S�� G�ƺo�nt��ҍ�TL,�u���ޕ2�t���� ��V�������B�fe&�����ҎN�v"5vd��XLJ��e�.$@ɐ��>Wg�d��8��i���]`�E���}f�}���t�v�y����n.I���>�2���4�]����B�ј�w*�!���\���R�@X���C�ԯ�xe�M���:{4̠Q��U��<�2 e�6�ߥ�c`7�֙Ԃ�LC��R�7����0}`�W�h�NK3,��"k��$����,���M�t}�ܘ�M�I#ń�{&aH�h2�CY�C*e6�d��
R��&I<��U����^bʰ#<F"����{�H�^g�����+�|�wt�&)�E�h�#I��v��B��vw���, �?��	� @�@P(6�tC�I6�M��)�U�3��qݞ�����ʬʪ���ow�2#�7�y�c����
<�M24�?�J�,`)�P�-���3^%���-�f��tU�5��-P�\���}ƕ�Jp'#E$�g�9��umY;|29��x�"�mզڣY���I�����2�=��+U����e�˻e͑�7���O�6�	��ؚ��m������Q�%����|����������ވ�n7"�z����Q�?�8
�ۿ�.�i��a�(��X�]��O���l�w?�߻G=�A~i�Q+�N���K�`g���5	���U*%�Au+�^Ћ	%(��^�رj4B)�wM�0�V9����k�X;��|�r�:9æ��M!c%KI7Lտ;��C��p�Vu�ņo^*83/� ����%�!(L"i"��Z�x��Pr�Q�9hʸ���y�K�Jf2���-G�o�3'�q@Em�H����EY�SF\�QPi�n(����㈱�eJb���:z ܅� r
�`��CF�+����BRio��!tM�ɲ괸^ ���� �*��BL��E�WU�W�v~���0�I��q�qS+q`��h��V|����7�-ܮ��0�x=>������A��o'�?="�������e�����l6EG�z������K/^��������Z��.^<��X_���P�^&��ܽ\
�e]��@��Ȥi2k�V|��"�H�n�����!��"U�����K�8b���Qo���F�Ճ*�)]M�d v��<�Y�K@�TK�N
�?Q�.�V�ɍ���}�w��$��^G�Pq
#���rE�������D��@zp��1�\�l��+�keon N��J���R�);�� {�)��l�RlH
����L@^W
��[�E�:��~�E2�F�qJ���}���tM�?�nQ�$-�ʌ�F�� s����2��u�5�]�.&;OpHs�m@�!S�E7��Lg�L��2�׎
�;��
zo}�w>�L����t���g�]s��q2[��w��j	��
�p��|�������e���Q����c֪߫���/_�Y��Ҝ�$%����;� ��h8Hze��@��P��F�Ix@H�"�5vV<��@UQ�Zf�;*�(�B��l��F�����\��z6���&��@^��:��-�Q�E&�8��"���Ç��1\I���%z��O��0�Gl �BX.5��ȱ���2�1.���3�Q!1�����H �E�Cc��V��~��~���'�b2YCy1�G�f	9�g�~����l�_RH�2د#
�iP ����r��X�DR;�k��u�룧n�B�Ħ��&� ��Ц�2{��X�������9��d��ɗ�F�fl�f�O
FM�Q��F�T���?�!��=��?�3rк���(k ~aaA���7�X�@�������o��ur\��%�3Q�_�ի�~*bf�{=��"ɋ$���ሒ��'�<�퍄f��
#-�!O�����xY�VP?���T�}2���`�po������\rʕ�'�Ww%���^������4�XKm��|��Yd>f :���m@���[���ÂZ�'Z�4��e;��K� N66A(�F�h �=iT��5��S��T˼�.��Lm�F�r5���E���d<�)b���F=�1!�H�0s� 4=�]H���d�� +4�ǵ�+�&e��n]$$3h�|�0C8�iG��Ѣ�t�J��ͺ)0�̉�{;|�D��8�����+F��LN���4�7o�A/��T$1�����������A�� �N6PG7�~7�~�#ԭ�Iw�tN�Qf�X�N��0��̈��`��
ş_�e_�Ϗ$g`�u ߨ��/����>�,Z����u�:e��P.M0��4�(�H��VI\6�n���uS�Ri���v�C�;�)����O���H�P��f�麙˳��X��)��s��f{W��!�{,�GR�/#��1��š�����y�W���3w����9ѻ)F�)��%>�:�՚��2T�2���1��?���TB��Q$c�׵��m�kW�U����*�Eu��Dy��5�������8d����^Q�}�D��Kj,�OntjDcF�����/����L7%�@F��B
�j\I$R��&��98��l2^/��E�EV�C3�X$�����G��v�^�BW~���TT��=���VǍ���S飬;=^o�{��o�3�1�য়��b=�۵L�
��k���$`��Uѓ������V�ݾ��)?ގ} ����T��U�/�_��7��l1{O��^9ȩ����������1*蘰թ��d�Z�P0phm�+J�ȬCAX�a�莘�6*�F�������p���۔����I\�j�B��`h)���h�K�L�����V�h�H�_�o?�I��� �^h_�'\Њ��&��~���x@2�H�<W��F^"�V��4OV=|�%� U�^�vW�#�Z��*�:hG)���U9_\<V����üB�b��}^���>1{y��/.=H�+�M����P������yV�2#(�1�M X�X���Z���l�Q`V"��)
���s���k]%��e#���fO��������@�����x�����5}<�go���M���Hsssc_<�e��J��%ƴ�/|��4���Em���?�z��
0�q�����=@;�W�!4�]m�b���+��ǉ0r�H���-#�r��R�w7jP4H/��k�(4���5t��-S��f��xm�*��;��A����,��,I���!�(���BB�����J�wM�N����"k`�)��1�#�����ۑ#E@�Q6�.�:(�
� e*��0=9�͆�פ�*J��e��ƽ<�I���� ld��:A -� ��˒(O�"/�AO;\S ��'o�՗�ގ��	�-K�,Wt�a7W�b�'9>���T���o�`l|q5�̙�oD/գT�LWȇ�7�%��팛��7no�U��Q֛���\7 �P�����M��wK,cȯ,5�[;����Fs�!��@�a��H��`����
`��	���e�U�B��J� .�;��"�D� �y�� �>1�׫��H�pg�¦J���V�V�1^{���)S�i����.��~�E��R{k��R�
�K��,��E@�UO�qEr�e>M�E_=��^�Vp�:��rn=��EƳ���6��5(�T5��.����B���U#r��@�|���
o9ŀA:S���`�.��Ԥ�C���\�\��4����ݻl��v4�9��Zc���Йf0��-�4�O3֙,��t7����=�}����n�c���F�c�ar����h�:`�`����n��]���c�^ȿ��?��m�wg���Ow�=Cۻ�3�Fn��3�DX:p3,96Y�Ĉzш"f�^8�Ĺ'���#���^/I�%|�?�F=�2�h�%��\�J�|��m��TI��ȀN�L��$"�ʧ��H�	SŁ�K��z��So�MQwH�a*�*#�G����l� ��j�����~_�̶�wh�5'�>y�Sy>���@��Qh���k;Cqs���exqP-�����gh�U7���!��kC�2�P��L[%=i�j���sg�q=l]�k5���*��u���&SY�DPHC&�X�[68�ߘ��l��|;"=6w/�E�G�n���0n#�f4H������!n5��f�'w��D~�{�Ό�;��S�u��>wo��@�0�g0�gff&��0����q�-�} _
���'���K����57�tum��$��Yf�ͪ#RÎ�)�4�
o�u���-��l ]���Xd�;O;;}f�-�_���Z=f?���
=Z���C	�� `�^gI.��R5	+!LѤ9J.xFVΠ0E= x�?�G��0� �΀�A�8��T�í�,i�`ø��S��N$�
U�8�$����S.��+Q�kD� ��B����	��Ir/��|��2�(l1?2���"��/U��[�טK�ܝ��ka���+�Nu��|���)�G���Y�Vm{��)��`�
��-r� a�7���z����#�[��lpϠs#i�y�%7^�+lsr�[3k���owLO�+@9���;���v����f�Χ��l��� Of��3 ?;;+.�?v W����y$y�ɱ�?�3?w�?���-�6�Rf��Yc0[�x�E?��ר�8�_�#=Ys�5�$bD+KK��T�y�L�8�)��?���E�0�hK�j�U_v� @[� �����"#�k�~����+0��T���i,��Iiz%|�(���&D�;����	2¡ *䇑�R�K.��^��rϷ��g4Q�
H�|��(��sǴ���&�;��˴F�;嘤_n*��V���lӖ8[7�Sh��0d3{+�:�?���se<�t2e��u�`�#�$���k+A�,�dc�8g��LRU�U�G5��$En�}���/���	<s�/��� ���fY�:��)��q'��s���I��C��v�B�$�9��f�O�j���9�} ������yՆ���ْ4iv�N4���w�
�K���[w�ܰ�D��[�0�t�K�aBn&L��
����	�qP��ua�>o/����몽X�>�
�NGţ�,�3�X_jz(
�GC�~l R5r0� ��k�Q��Z�A#6��P���*�13W4�{{�N\B����#)��@�Q����� �W��P��1�Q"���0�� �j"Bd��ĸh~���[O�0K��BV��y���&�<(`ϙ�U�wT?�	c��d�reV'Ɲ�t�7^�z��R�d�m�ϵr ��ׄ�f-�
�E&)�H;ʐ��L�p�]�2�޷��Gi����7�=���ͪ$o��rr���Q9J1�d�����Q�?,��F��s���q�󳊕�![ {�9�)*a����<���zd��ɱ�'�/�����s�<��s\��
z聓��Pb�0��a�
Ck��l�ii�%:)�(���ra�~�H�G�l�[T�BG�U��(�P<��O.���ʥ��.��t��YD��X��>s�D%�1�n{T�"��,Z���9�$�H�L�H�3`����H�T��a��.�J�..M�N��Rf��l���ZD��.�ԛԜoH~��N�-�
ەʑ�2R!�&�K>�Y�h! �Ǎ��ΐ�%�j�G�R��'�+C��
�D� ���r!���1˓�βe���U��V�-��Ք� ������5��C��HH8*��b���7�y�?s��L*������m"�?�Y ���V���^��187�fy�ǭ���h���ip��\���n���*Mf�h�J#��5|�G���8�ןx��6Nq?�ǃN���O6�/f?���̰�Ξ*Q6l���%Q����2���ئ��Ye5�ű�je�����t�� aI�	4YFZ��䮤^�ҊO�"��Ow���� ���*���IJ���Y="o���l0��Iek���9(iK�,�~�.�40ZBu�3p#��.��L��)��yg��9jo��<1[4H�k5�
%�D\�jI�:� (L?ְR�FI�4 GF�F�M��`�FSF��M��}�L\�۩n��̔��Dd�1�S[A�+4/��� �4���Io/x+AT.#_��jb�#@~=����/�6�v�F��xi��,�v�a��}w���@�zǍ�$���'??H�`��~#�p�}�u��ͶA�+cW����ɘuKR�c�W+y�$��+���եSђ��]£0`���Q��K/=��ꮼ����8��e�@&:([n��f�֮�����bҰ��|qhV#��3�l�ԥ*����A��D;-eZi* �O�Z�6A�S�%��)7���Q �G��"���]4��T�R ��2a ���P{1V��i������R�6C.˕j�˸"��� '�^!���kb}�p"������_�ڔ�BR#�yg
܎�^\[��b�Vu�8H�v]�~�gl�d�ءA��_d�����ڭ�jΛ��V��� �8�\s�st�����cF$j��g#u;ɜ�i����w�8��~3��N��g��B*�A�����e���=����Z��4=Ͽߒ������g� �.��`��s�^���}�̖G��ڛZ��\@s&!H�7���,���q�.�U��2r����ǐ").�ye@����Iܧ���
�7��!8l�7�#��x�B9*>���˂]G��F��<�$c&�VM.rf�M���;PwN:�(��L��`���M�?��>�2O)�u/7�./��-�<�;
�$�j:/�羧���e���g
7�J��,�׊]��*Ta��rru�1�ޓ�n�<^����p&V�J��H����2��'9ġt�r��f3�AΌ�*���`���H�,��Κ�����M�mc|of{'Ǎ\o�qн8jL�fES�[eٻk�/R)}������6�~wMo0*��v��s;O_�8y��:�XiQ�>`0v��V+-~��""���{)F�;�k��0 ���4�*`Fc]��f��(�LsB,}b��Y�4bv��"�$0�2��^I�	rչI�L�[=��"���Q�8� ���4�����uFAJk!ľ��G]{w�� �H�,W[���Dkkk��s:�l�jH)�݁�4Wi ,�6�
���Z�,. ��?��T'�$M�-��ؑv(}Q��q<������g�pͶ�k�'�5Ȗi��������<����33.�l �*_a��������䘽���B.b/�lZ��YGS�P4֟���M��I�w⸝i�$��ƻ�;�כ�t�q+u�ˍ�s'�?j�u�3+u<�l�m���>�������[N��c�@Y�N�&e� ^�%�hч��^J�����GQ�S��hHOW�)����m��sTB�l�ba*Y(�0�T��D�&h��	ݔQ�3 �4�Fu�:�k<٦\�L���/"��V�;]>^u�����#ĳ�Y�բ�	 r
��z�8��_���qk��P�C�o��QD^��%��88�B����/�⇒
*."���,����DyI�+^NB�뮑��q}4-6ZYk\;Dc��L�t�UUp��CV��k=F��or���>W[���EQ�y�4kH��L5���Ѵ>����j0٢����� ��u�I�~�����?+ǭ�s�ŭs�u���vY�̓wߡ�	g���v~�/߅|����vf����溯��M4�"0g���Ր;�Ra�pMHWa߅ho8��������̀c�7t�k5�n�g�J}�{"!  .DJEs�E�����R\����� Fe�ĪC�����5k�q>8R��>_���:��<Y΃!� h����L�~F���h�����&�lG���c|R�d�G��z�P��֑�權�2aWa� G�),RD^͸O
�c+n�B��蝽�X�i�"L�O���= /�_��,�`�����h}�4��uWXa��J�r����|?�$MNC�k�!s��=s�L~~T`�Q �<��o&Ԙ�Q�c��Ooc:#'g��J�{��b���>�я:����J�3���~���������lk�����4�R����5̊���L��x˓��-dP2���8���z�V��AN`yK�S�T�̐锼̹SZYj��U��=���]qҠB/L��*hVj����P|�FCW���h�����Yc K��>���v;�- ;���l��U�:�vo����2K�;�IJuc����S}!��Ѥ�����U�_X�����j��c��QH�Z���'�P��(���	D�:;����E���#.�F�K���r�<�5�@�3�B#e�{�9����3�=w�c�R� �²q��®%g����q�e.�N(Dw�$�]�d.����$�3��Ul���@ϧ�88�D�c����y&_�ɗ�f�(o�8ȏ��n����Ĺ�F��<�i�|����f۴��7�=6ˁ )@ֿ?賃�1It�Nz%{�>a���������n�o�a�NO�����'{+++�O�6�v�C����(�,J�pG���`��$A��٦�ّ��TC DMG�4���^�0$���� �:��.]�m�X�f2U��O� a�-Z)���4?{J+�!���H�� � ��Ǫ����iB	���������P�קZ5��km�x~�3��M��G=z�b�n�嫫��~�N�<@s��3p�A�i�|��+��IF��Q��ۑV��@�#�f�q�Ŋ{i:�M�L+=�(�uдJ	�"}ݸW$=��i�uؗKZ�Z��Xਦ����B5}Յ εy��<w;+Gk!��K�Y��c��F�mu`n��_�R�׃^��3���5	�o���N��uS�]Ɲ<���Q��'5��>���_)7�|��w�1�:�__���wj���|,~���
|ץRE*?�4C{��Zl�kp-3"]IR0�1Xv����
1Ч�����K��/Y.��.c�xH�����3��ÃQ�+ȇ�:����T/� ����#Ɨ� �����Xt摱r0Gr:\u{��P��8��s�C�66is#���R���is{��c�_�X ���xO+'��Ty��~*e��z�C�Е���5��.�L�B��^��̤2�d��
�cU^f�1��\�,VJ@���1!Yݝ�ckG(0l�Y0��B��RqlOI���jS��)�n��|lX�.g�Ke�_����������$xM�a��ފ�F�� ��̾��z3@�F~�f���f����nu��ѦQb��目Q�}�����vw�����---�����#��!��H0�o ��ѳ�]�p�fYG��t����^(j�)^"9�.�z��d�Z��ʆ����]�a〴<8`��T�F���֣��Z+h�Ki}wD=���mvb!���G�f�f��e|^)�cr���?U��aq�=��=��sߔ�+�A�ϾRK��KT)�43W�8ۦW_y��:�>z��G�ʕ�����S"�R�����l�9U���B�n���67�([7�X�q1�wdb+^�+�LN���,��kǨ�;���g$���Z
YN�mr��45��Y��m��"(G�S�r�)��:�٠���s��1��/鯴���˼]��[qG線)��{������2v9��\8���lbػu�Ln _���k׮�9wMݍ�h8�n6O��f�)t���L�kՆ0;��Q��9�4�����\l�B;p�X���sN!nt�u�j��u�9��9�z���ܩ�w#ʢ�Y��|Fo���W��3d@΋���-:��#xȇI'W�t�3�,��Y���k��T]jI�'T1�	�;�2CՊ/*��ʬ�씫u�52�y�~�ڽ�J�
]Zݡ�����u�z�*}��eg�W�p�����_��.\2�����H�2e����8��NLn�4'�2i׀�ޓb �1�I�Q�����?}�
u��c4����Q������=��/m�R{Ǡ˨��u�=cQ�I��;�I����|�o�8�{X��V�A��0��;q�]��V�krpX�ԭ~6}�����AFK��!=p��-��@�N�bx�ګ�k��(z�Vd5з5Ս�N+�;D%�s^a̴>�t��y�fǹ@n���5_����]�l����,���<�2��ꋼ�G����fˋt��穳�b=���%��_��X~�Rf��8�u���9j֪�i����uմ��Y�<C�E����r'O��N�"����k�RB��(��^�L�6w�9�v{D��'��$}���N�qz��.E1_�ꔉ b�ǆf�8o��G,��a�P��
x����doU�G���ə+!���¤�Z�����V��M?44��dr�j8���0�1��՝�F�� ����%�ևxt���&�� ��˺�&��ֽf���L����T�_��2�7��r'�A�v��|��6�w&p� �Q�}�g"�Y-��p%qP�c�v�v�0Qv666�_���?���wgV�����/2��iwgK�j�%�)�^��U�Mf�Ȯ��iP�JG�
�b}W�k_,�J�*Uf��m�Y�3���ReY����	=�zէ�K�����ݸJ����2[8�T�����[��W���e�)l�^�M��y�'g�s�y6��v��?���}N�V�Lڻ����zS����B �k��k�����5�*��&�?ߧF�yz�C�]w���k/��FD(Xƹ 2j�Q�2��C13@[-��d���Cu�EK���4�FR(s���T%3�������b�>Q�ܴ.��^�*l4����pZn�����ZG�70L�0����*$��4m�m�<�e��>&?���q�%&3mPzjٷb����v��N���q���9�r����c����n�'��9ǭT*w�1�Iҋ�Q�j4(pEr`�vE*����#}����씺��x�xHf�q��2�T�5�����<��|��^��KKAh���������|�NͰ���2Z��ҥK9%Y$�rla��Y[�&���^)QeԚo��{1�W���9"�Ct��������5���ymR�F"e_�Ix�g��t�Iۈ�uf�]z���t����裏ҰS�����R�#)���C�,\��U��cP�q�5�l��c\6>�v�
�i�V���i�ZXà��ҽ��i&dP��恊�ƻV'{�Q���7�M�]�h�%R}��� *�p�S����g�Ŭl4�M+�Հ�ӻe䪙|�ov�o5���;��z#Ǜ1��ٰ�>Ihl���N�>���}�E��i����@��V�dy���U��v��RR�:۬��4h�k⏇?�T���������G�z���Ez�:=��O�I<Q�-i"�E�c�r�Ξ<� <���O���1��w��������R��m�0�hq�IǖO�:̀�n�~����M�^��Y��Ef�u>1/��Hr�+���S���:y�85���6�=�|V�-��x@k�v�|#a��P{ю)ϥN7�j�@d�s6llX\m�H�>�x(>zH/�`mLѓ#Y7|L&__��r�gc���=��;{�*R�!`���$l[\,���*� SW3e���t4T��Zi��<��|I��ڴ�U�9D�i������۾V�m�Cn�7���2O� w�w~����p�.ԭ�������2���EG�������};4��3=n���N7��cX��������;S�j�ng��';I�d�R����N�����w���E=v���=�*3�b��ϡ�y���Z%�i����U��X�� ��T��;� ]���Fb�8R����s3L�_ze��h�u�vBs�|!v������U�J/�8F��&uzm>d�4����}���m��]eC�*�r���T:^���(j��O.��rX��8Kq�����	ya*��VIG.]xm�._ؤ���d��&�0�L$�F�D�^�!�� �� �����7�U:4M1q�t(7�Kr��C4�d.�� o��z� �횵����bџ�a�&��aܤ�$rVQ���Ɨo�w�(T�g����M`/��,"4�9��������e�L���}7����Q3{��;333�O����>{[�5�|9�f�鱹si藼$�����դ�l�^�h��:5Y�*��x��	:��\~�̠�H�$�x1j�2Z:6O�N��+�.���z��
|�e��o���hww�P73�[]ߤt��FgDI��&��}~�Ì��v�^����t�饗7iwg�� �P�W^}��\�F��q�d��O5(��d��D+e���������!�y�Q��y�[���y�J$5����3���C�ƐJ
ˍu�4+U��X�m">�ч6�A���J�S@���X��xٿ'���W�F�k^���fo�ž�ǌ��dRh�,���Q��� n�������{O3kx������M� ����>����v���3o�8(��Fc2!bzv]�/���̙3w�]Ô}O�(d�G���\IGL��_Bug�WEXf�/TyYf��0ق0(�m0ho,�R:qr��ZM�������b�#ʨ���m�]b`M�r�D����mv�7Hh��W>G�$[�g�;T=^���:��ʅu�r~��8>G�3U�Ӯt�
�J��:=�`��6�bh���(�+W�����X0Y7��_P�N(�Q�2����v�{������;Á�.P|�Je�'XS�L})H29�����<V`r��{Y��~/:͂��_~#�ސ���c$��<3 ��yҼw���mUx�ϡ����+�FFy°Xƾ��XF����1OgBL3���fo�};�����o�~�����<�	�a�J�?���u״�57I.v �(�]�\w�ύ�ɗL�{4��,i�+T�!E�>b��{��F:%g�>�L�AgN�hا��	{��S��˫�1x�ϔғZ�ei�g%�Q��a���-�b�ZoK��� B��m��%j̵D�fwg�:[Cz���D��;Kg�̲!٥!2vx6jT�c-�|:��ia���2}�{��s��'HP�*$A`w�P�͇���|�D�AJh-M}TC_�l�d$�	�<�D�Q◅d�{=W�}l^��=��'O�JY#�<^�Q�0w�w4�ņ=�c��U�Zf�L�O��y�f$��~e����L��|���T�zBD׃�ط3�\��(�c��=�c�Ipߩ����;9����L�~�1�I�պ�L��W^L~�Ï]�L�6��'Q�@�y��F�����Ï�C+��R��ez���ڕUI����x�O���7���hc�tm�{��_�4H's�OrY�އN�?�A�2����������� �"iց̼A'��[�{�Y�J%�Aw�N�,��ph���ܡ���fh8�PRt�՜%�O�`��}�D���^x�=��K��C�� �� 
.�RJ�l�!����o���%��w~̬���fо/cw!ЖHX�,pI��l��R(���J[�6�.��˞��la �d�\���ڡ��[��@�5��jd<5F>Aν��+Uxp7eb�\�UP�!������5D�Q4i@r�?���Ǿ���}�6��r��V3�7����yo���v���r�\�=n��w6��c4�"�+�3���@�;��=�EJ�u]-Tk�-y�B5qȌx���L;"%�`6�ʅ�{�*�r}�`eZ����ڀN�8A�C�Fmj4�����љ�T睍����]#�Hѐ��xD�@&���w�"-.�c|F\?ѰM>� 0;�u��t�x�ƌ�8��3�34���KW���~x������<�\�b��\���l*N<+!�_jн�����<=��,�$U���J����Qj��	�4AۥC�e���{a]ĝUB`���Ƃj�13�L�V�ʬ�����ˬ+h�9I�?u�2���QิG��X��+�H,>�����9��v�-���Ŏ��m�f���x�o6�QfΤ~�A���J�B��v��@��{˥ ��*�L�y�ߠ�Ff���~J��P�J��䐚59�#0�(So�lnv)���y�l�`�S�ՠ�-��]H�v�m\iS�����e���qWhm�����3u
K%i`��q�*ի���$Sx�~�v� �f�t���]!�ܢ�Ŗ�.zxUC7'�����'��mB�vq�B��Fh�Lk�U�
�<po+ȟ<9O�N/�_����J�b�F�R ��Lc�hl����Y5���սarK��t��<��I�^m��Bst\aM���KU��9�؎ޛ�X����V}ɠRT��?WfUp?!^�=�]_3s
W��B^Bֵ�]�J�63�4�gB��>���T�}���a2��)�{������ƴ+�f�b`y&WE�����ٟu�������} �ol��y��4j��8�H58��!��)�A0�[�
�c�`�,<�Z�NP҉�<�7���ac{�����(���=���?>%q �^E�%Ҳ0��0���؈Jh�Z��з��?x���iqn�6ַ	]� � �4�22�23�^o��y�ԃ���<��� S�N�:��ȣ>��3+�Twiwk�\���^D��}�Yz�4���gu�:�=�'<���Ld�n����/���H�[�o;Gg(_U<]�7pR#d�+Ы�[�y�D��J����ڀ�c�I��F�X4�%@k��'�z�q�r�26bvK ��v��؉P�����{��EǕ�td/�(�xF���d�@�^��/&����i���U�G]4�6��́�_P]�b�Z�.���6\Ww��#�3v���o�U2m���
S&gp��Ȥ��6%� �4eNDR��%L����T���|j��i�7)�4����d���Z���k0�;�~����m��y���8��C$�t��F�e��Gg�]V�^�@�`,��3�������A�ۡ��̽r�ʝu�t{;N:�N.�+�*�e�6A����J�8��+�� �v�'e�x!�d�7\����]�S�/x���/ef�RF� #���<&`ǭV�<��.::�Q�Se���?�r�Ά�G;�tm5��;�Ta#T��E6��cT&���
�!��,�w���lTx&��فG��10�̈��� b6*�hf��U�sg���96]��ܤ�����������h�"��D�\(*­�"$xP2�
�H���k:�B�+g��E�^*������1�e����Q�v}d���L
��6�V�����V�x�bAW }��À��<nY����$� ��SP�%ƃ�  ��$�0��闋�q�l�u�U����;��ۓm�&���h�'�.���댇�*��7{<6�_�6���So"r�8�x���eu�����~v�ɘ�a�}�cy����F�V[��Q��[~2S@cZ�1����7�����q�������~B�9�J�'���
��LF��$E.yW��.�܊��ORi��xe���b%]yإ� �=&4�Ց�P�o�Q�fg�꧚bA�pE!_~{�#��H�,��H%8N�Wf�R�l/��S�t��qf�[�U*7f����0=���&yi��W���w�~u�g��P��~�i`�j�i���}��,}���[��Ox?�t��:�]\�T�X��$u�;cv	Yת�#G~B~�����v8�8�r/=�|%Y2��C��se#�*ῥ�ա�6
����A�cj`�A�mA��#�"oϕ�M ���y`7��`�<SA{F�İ>��� ǵ�bd�n�3���>zz���x��>����E���(��?���.!���h�{L0|�j� ���y:��*ɍ�j{L�6e�3��b��yZ��Ifh���A�m�GxO�e����yE�S���1��Y���M1&�Hn�x�cTp��=������������s�ׁ��!�O�۠z��L�w���Vj����/#��@�Wnj13M�W��J�t�k���
IA��AU$�9�ZUm ���T�8u�4����%*m�k/��M�� c.		=y�5�������/�_�sw��3�3�Yf��4��է�;G�fF�~L^�ĳ	��V��ɨ+Z<È�H5x���5�r�IK��A��v���m@����t��WT�v��2y�A�S!Cg��hը_��fas㛾����*��׹��_ǙbdcA���"��'�ˍ��1
�^�[�kgm�fif�Lt����ˣ,����1�f8ZIU�&�`���I�j+u��'�c��E�`�k�m[`�g؟ݧe��Q�cr?��)W��r�F�N��{X
e�j8G|f{3�{)�/Ȇ1mX��xzfw�L#<��?�4=��6��Fؘ�֖�O��k3}M&��u�H=P�g��6�jH'	4k�>T��;�B���vg�W눪m�p�.�L��;��(��@[�<�� �X�#+1 ��O�h\)�$BXsQi���ϽVR�YrCb�m�p �(D�x�C}��UZZhQ��s��&S��H�An�7���i��I�te�^�p�N���x����x��J���*>pBW*�WؠP�8��F4�R�ңN�]Y�B+K���I��[2�X^���pG��;[��k�1�_��+[��#�tNJ��$Sޛ9��HL!�bn!���Ix�M�%Ȫ����}b:H�m�K���5�?E�� ۂ��Uo���e�L��!5!��2��@l�Fऒ�{�(�ib2��r��}���d��_@�T\��ρ�O����-M�q��Nu}��+��}i��Z���`zd��ce]vV0�J�4(v�5]i;��f���j�a ����� ���˹�1(;ĳ�b���o���[��e���z{nv9{?&�e�����4Ƚ��&��sVE%�^��̸,%�����3��Ր4)�+�cإ'}��}��f�7�ɻ������/�qP�o����(�(Ni��YZ�_`f�JaO���`h�Tk��]Z��)|�?�HaD)?h�=K!3�LS�H���3c��	 �j!o+�����Z�ev\�}Th0�)G�6�^tȬ��"j�̲��3)��/]�ܫѧ?��t��(�̐S�I����9̦|~y�H\
	aP���c������K��Cϑ�_{g��fNS�3�k�#�m^�����%��E\���9��L�҈U&Y:�^�3�t,xE��ş��>�5s��-��47߱�:���ar�GF���u�4(@��&!�;����wh܍��x�K���Q����K� ߣ�"�J`.!O��� ˜T��@έV��g2=# .�/�������+��Ƅ�'/�	��� "�U&U����&��Vj`��ˡ׀���5�X�F�{���a}��Sn������F�>��4�?ȸL3��ޠ�m&����ǘv�L��n6�j�Tc4��=n<~>�a�����:y����y�;m��3�i��ј�����t�j~�_��ׁ|��wK�Q�)��P��	O9�A�To-��{k<E��/�a�T�b�k-��˂�hfݔi�ߗb'4�.\ts����4X6ʤ/*@�V/f$�fժK��e�+�N/䗨�L�Zp��1��@?�sm�C�N�K���Ԝ?�S�%6�(�ʥ��(BʙQ!����t��A�g	a5`��/}��x��b��������g����0w��ȡ��U�b��vG�  ����,g-N�|���L�pG0��bB���坉[�d�1��)LO�l���p�ˤ02��Y�]��ۉ�Bc�W�0��QAg֝{2[|���
a8�,�+1l�a���ĳ,�Y�m����h��H�-��/�eZP�ũ�h@*7���|��J��ά'�lnl�u��[(���6�'Rj-H��t&�?�����aܞ/�F7�h���kM1����|�9Ï�^T|n�d x�o>	�����?qmUcH�>o���Y��y�e�B�.����Ę4V��Ե�	�A3!���H�F�E�A�dd�]������}��t����Æ��l6�\g��$���ͅ�@��/�_�E+���_��_��l�j5��}j9�Ж�y�����n�P{k��~ Λng[dz�^X�ܥ��R\�US���g����6#�1�g._�rN�"�|zd�X7��@*���_�!3�}?�:������iĠ��˝�!�A�CQ�D!�' ���
23K�ŕ���稊kɳ�:d3�<�l��5�B�y��vJ'V������)�5���x�XMh�UА�OO���ԙy�rm���u�����T�5�z������]���~�L��d�Hw.�%&�.-�Bj�f��O瀞���6$2l�P ��3�	O���3(����V�.��}6����te?�RY�m�h4�\a���Lڲ_�� ���w�]Y�cX��]�m�s�m�����?�;���p]Y5���(�և<���2}Fh����i�,�x��c]��Ђ�u=M�P&�99&;gYw��	��m����Z�xZS�{>���w���#ȣ���y�.<�����z1i�j�\{�_�ۚ�v܊ќ�����5��$�v�ܫA���sZ*�8��A����~WN�kR4��*���*��ʵ�f��f���/�����>��7)(3��:��t�S��(��A�Ā4�h�)D¸?�3f�yS�1�
 �PĬKG(
�lxf����S�"�4_�*�~i|��oVY�A��a��wwv�e`��!�*�0y�:Z����	 �����Whey�N����4�N�_諻V`��)���&ȌT��^�K�i�.w-���4~���H~�i��q���T��_h�7M��-R���;�nбcs�;c�v��-W�Uy@�]����}��	�� !Qe�F=	 ;���3-�_��m��9���W.S���@:�&Xw���"A�S �PN�l#HX��L
�5������@qm�����:mllJG2�ʱ<�Ë�[k6��`�]�_���mYfiqA���}�C���];c�/7����󋼯�|W">� �����������6=��bx�����,�Q���J���-c��5�qaaN�X�����}�#u�9���1�eqW��p_��{�.��{1>;|�9� ��f��ǌ{�g�k��ol��w��5��j�33u�]��k/�wl(F���5�ե'N�0R���\S������=µ��5��t:cck�e2��^8��d���9��t'wf����f�����-�;%fd�*�����@hE\9��]� �4b��"���{�)g���"��hإQ�e�ҧA:��g}�� -�٘��t����iT��<O}��>&���I�N=H+�ȟ;��Wb��۠� V֌�=譔`y���q�9����M�vTt�ŗ��ۦ��:��ǉ0P��8i����^���^$�����X ˤ~�����[�R�A!��G�g4�4��n��$�P7���&��OL?]G Rض����S�U�G!���ȕ�h���װ&FP��ſ���ϳ��"���3��(��$c��������Θ�!��̑����Ҳ�Alo�2(������������?�����t�_8M��Y#	0�̪����5^�k���GKKry._�LO=�������\O�< �C�sqqA�!^Z,��/�-Ly�W�Μ9#/<^�J�* �n���ŋf�pߘ�bF74l�� N|�s���X/+*�q@p�<����m��W�B�?��S�`��ަ?��?�D^` ���@����q��+a��|b�Z��H��'?�	_�k���}l�`�'��U��ll���� �;��Z�wʰ./�;+µ�盛����,���S�����\�e&t��=y��b�k[���[����xO�.\�Hw�uZ��1�ӟ>ǟ�%���W��w2��1��������L�={�����Y	�j�/�5�N�& b�$�{�I�_����U�'U��Z@.p,�U�4������@}f��6�F �.� �a��&|3_�}�@�0W�B�x;AX�N�H�� �R�3���S4�t7-�~����<���gV����	��)6hs�(#��{����S����2H@ ��,��&�#�Pb&�ּ����ª<����м�5��C@�
��6h�lГ��R�X�æ�~)&����'��>���_r&����A�&��J_{�
kNK��h~aFd�/�_v�r�%5#�~�ׇ�g�3��~�*]��%�|�"]}e��x�e:~���z��Z�zU��XE	��>����I
3�U�}+1	x������g�ۥ����>�:w��Ua�z��K�������~P^���WD����?���_��\��_~��{?}���]`�1�����N�<��?'�MZ�`����|�~�����O}�>����-�u����/��������0��Ǐ�AxY������%�y���.F=I�m=�������3��<�
�j2S������o[����W_��:��o���	���J�_�}���A���{�����{�x�$�y�MPw���wvvLp�?��O���}��|_�eyucm�s�='�O��O�Qᜰ��49�I����u܇����5���}��zum������tZ���NWf�x>1�}�	!��ҒdG�c��J�VVVD*������>�.�����8�\W�D�x�ow\��{���yN5 ؄v�A0`O�Bc2]D�^Q��3�`����[B03U�C�ĄA�-jc��93��G����g��u��I�{��v$�0�*���m�x��yZ�]���*}P[b@��ā�V��	!�o���\�Ir>�p�f� �~�!�X�|���~���5!sP�#	p|#@�ۼNveU|�Z�6����$ē�I��y�L����l�/ѦSd@Ϝ�gd��ێ��:aC�u���}��=�_�1��S�Z�?�C�>Kj`٧��ۥ����ب��g���V������3[t�5�O|�_6�[�=�t��u#���͵(�k<���̤��Z���5f�k���t��k4Ӛc��!}�3��"L�}��~�;ߣ�gлt��8/�c�=Fǎg�`�s �?�a��7���^������t0�=]�?��?{衇�;,��پ80$��������(������	�������x�O�fcЃQ���:�����o~���3���x��
�� ���4y�������w1��|��_�cp?u���o�� �}�w��tr��@��P����#���p����<��mll�T��[�y���#lv��_8<�Hx����|w�����A���o�~�z���W~�W�~>�/��N�>-���o��o	9H�D�	>����~ZfH����57���d�|�.߫`mm����͊�9qP.��k#��p�Ճ=�s��sEn���5��0�ã���?��)�w`�v�)1R0����쏷٨�6�y�ټ@� �x:C���1{kǨ�Z���}��e���GY��=H���O$�'�V�J����~�ϴ/U���{��Y��lY���$u3�ͭ�"ߔ�T��y"Y3�A|w�/������҄n� H�L���g
�0��i���!75�'�{6��0�����<�ݚ�E��-�j��,��:l'�}��p�TE~�GO�Lć+ha�g=%�ڝ!�Zj5����&u�a��y�O�3����D���`�	mu{��|����䧈��倬@�5p�Ao6��L(K�8��Y�k^�o~�[���g?�L������8���X/�� ���^�'V���?�� ;��׿�L ��c��˄����u���ܹ�%'A�Vk��i�w���y챏ȋ}���ϣ2 �{aS=�i 37� �����ws�r<�?����0(脆���h|���+}�#�k���#������G��G?�Q9^�>\*���Q�4?>����l��lu�]�rE@��X�,�ܦ�� J�1F�/H~'�l&g'8\sK"���D�_��\_ܧ�|�#�`�/�����?�ʓ�����L�Ķ^~�U&��\�?��?�uq���<�ܳra`?���k�w��Dv��00l�|ڐ�:ߗ����@>ڍ��(�����^�w�)��d���$�d�EA�2��(�6w�jh�K�TH5s��[А�!�J��������Ǩ<�BQ���;�Pt���f�2�3J�켽���#�mA���^��97:�����1���X�+���-ș�7D�Q�NP��"�J��ZW�I�?�����"����iB
�w3G�2�W�8{B��5~OAr�g��Lܓ���k��a����Y�6Ks$Ek�Ȍ�+eHCϲѫS�>K�
� 4����y��ݎt����}�>��*yu����҉3�2�(b�i�<�����cpm�
Q�sS*'������.�_�� ��K@R8/�g�K_�2=��������W�s��� 4�+\.?��3���/~^�`�������^$ 7��׃���|��ya�`Y���/�o��o�K��/}�����\�����/�_4��Ƌ7�3����ȵRq�q�?�^+�f_V����0 8_{�}�k_��<�]��[fp��X��~�CC��Y�� ��W�E1� �b���`k#0ĸr��� C���l
�㸰���>/ϥ5
�	ay�E��E<�1	<�4���>)9a��1������II@��i��o��xG�y���W X�pF��F�_}\��^���s�g��ӟ�4���������;��Ø.b���a.�d|��\1��.���(���^,�0zM�d��I�Fb �B"�qMfq�����`B�Ȫ�W���,����3��{TYH$�� <CI6+�=��Č�K�4�GS��3��Ld��w�e��>ٲㄗ�r�y��ؤ���S�h l>Fn'�~��j×����!	���L7�w��>r�?Pl�Y����H���M�FJ�3Y��*���'_Ȭ�ƽVSې[�nX��F� 3�$#iww�ʵ%3��� ���5��� ��JU�蔏!c`���՘ټ��}��g����顇�g�y����J-6x�~Z>5/L��!�Q�U�D�e���`?��c��}���"En ����[���P^��>�Q:{�  �?���/}�ߙ�^��vyy�~�WU�Apkk�-Si�V�i�"��T6}L����e����ߑ��z��ֶd������&��������F��5Z�[e�b,��������_���Sp���u�����������P��׿%����S��#������|~��^�W��>_~�e��5�V?���-�+�pm1���1}�[ߒk�{��{r��M��m!��}�������_��_�c=y�d�`�6���<&�Ku��i���k�]�&F�O�ab6��W�������?"1T����`<��Vh�gYpw�M�}�3;S qX[[c��W�����������+��,M������$�s ߜm�����t�$/��ƽ�z	R��'_��Q����i���{.���� �y��$��]5�?��Gg�F�!O��^La�M����"��`/)H�0c!���!f�j��S!�'��#�l���6��{�{�je�9��j���H!�H�qP�S�\��X�ܑ󍢣�ybPg�.�6 �n�ė	�8e��&�Tp�rt��2�O�B�����������D<O+W�b(�)8�j5���
i���5�,m��F���b<�uK�9�����! �����M�wLef����t�b;!��e��=dV�kU^` o�l<�T����9I��˃��K����/,���u�F<h�/�w��]Q<�u�a�[�����C��O<!�������7�;㓟�$2d&�!��zU�AP���q<���'�+/�lS
` �����5�����ʞdS���}�50sX~�CR�W=d]�c``yܛ���3�{B���/�u� hq�Hq��65�oF��`�x~�!�gf4������/�}�S��4J<#8�˗W�%�4�_��_�g�G|o��'ą<;ےk�Yb�+`6�裏
�O
���N��ۚ	�.��vm]\� \��p/�";�g	�}iIS^A���S�
�����e^�4}�3��g^�o|�kt��Ey�`l��v@������6L��u�iݹb�������eZ[_�2��I�H�:T�s�B&d�h5]!��qj���o�Q�V��ѮERx��b �J�X?�Qich�X<�
�<|dǄ�������.G�LTel�'��b����]��3o%�Q_36��&���-�w��^���0��g6��E�lms�|�
�VE�u�7�=�Q.����\����ZEg�5���ɇªL��$�=���ل�Y@�L���udd0���;�6�рmf�L}H��H�Kha~��jI���R�wy{�<C�H����!����>>����p�9��Z�ϙ����� {tby���'�5(f0��U&�vp�S��!K2��a�������U����JC�Oǘ�۬� G�Cvx���G��C��?�N	P���3�������������������Ut�����De���uĵ���� #@ܿ{�(���s�s�[9twuι[��J��d%��0��<`��1�Y�Y��b�0<�{`f��l�sd+�nI�Su康��4���w�v��3F�]*UWս���/���ߍe��n���C�f��̡�Ŗ!�i�c�(�[o�ՠ����C�q�(%ޏ`���/�Q�lܰل<Bghh�BT��q���gۻw�]'������Ey�գf�=zB>�_���5�_(:dttL���)�`��k��*�b7�BCi<�����~P��N�N��	��"!_��������7B�0
ϲn��yB�=�B=����;n�=w���ò��A� ?z���c�B)��@N�qQ�C-������*	mڼN��w��ߣ�b W^u�y�>����l��
#���?�{7�{���B��*�ztu\7u���$�˫e��r;�7��e�a��^=� Z�l���%I� :,��;$I��a'�N;eA��,n�
);	�xVC+k7��&ah(/�#'��j6�?��&��	��Ϟ���d~��-La~� O��͊���L5+M�w5�y�U���I�V�޷%�q�*WR��+rq��z��4;.��郐z8d��*��F=.w��ܒ,-�MP�&TH�dh,/�*ԛ���OX���s2�vLV����y=��RY�����+.��Ų��B[����|Q�U�w�Z����#��g>'�
��y��߬l޺Z�hv�b�� ��JPe�H��[�m��<���R-W�y�����栅6r=����*w�rB%�����w1���/��	5B�=X�.~�2����xFG��-����fs!�c���I�y��cFP�c�vٲu�	��\�'R�l���p���Q�����e߾}fА�@�ʿ�=�p
�Qչsg-q�{���k���X�n��޽��V�BՊ���²G0o߶�*��@��}�h�'<�#�52�o���-�D}�?x((sK��<��f�*�K�������>b�|^̡mt.�Y�S Ύ����B2���y����r�Bf�i	nܸ^n|�e�zaD7��N�0������_��S���������(X��dRl�:����{����<�쳯��SoƗJK���V�D�yBTIU��8���� �Ý�
�NHy+^��P�����8~����l�|CL�[�2�9�!H�ag/_��G�Q7�?1 �Z��)�L�K/<"3gd~�T����!�R��T��]�H*���&TK/L�c�["މ�����~������/[~��H�HV�.zd��˱C	���@U	���TC�}��L�[Pő2�'�^W\�C-�Q�Y7lf�,�/~�!ٺ}�,��+dl�J��� /I��HV=���^	zU��KS�a��,��/jr�E��%�Kh���*��ɴ��h�zpT.�uLBሻ���%)�y��G�S�����7��.w��	�W�[�Ѯ344a�b�z-���������gB�p��`��-IR+p�p`����F`s-��Ni,E�d\s'HיW�G@��G��vdt�	.�#S�X��铯�ba�*M�걬y~�y�z��#(A`��'~�����	��:۷�0�;1�P1��(���4%8�j�=���=;Ͳ{�\#����;l�jB;����VD�ƙ�P��'���뮓_��_5��<��-mNAx�[�>���)t�x��G¾��^`��γbt�.��UA��(@a~�3N�B���/}��x�8/����Cܞ�-!˻��(+���:>lD��+ ^�
z��{.�5k��O�z-���L��K��K�������շa�r�����}����cv�)��L���ww� a�x�+�w֒�"�Џ+	5>�(�q��:��6���#���/Ӄ�Z�veAΟyUf'����ڂ�M��&��.���Z(�E�Rk�B�i��@c����6⒲�)��S���G!I��AXų�c���]��Z�!�Ԉ|�s��ٗDrٺ�a���kxF��&�p~FΟ���RST����h���m��e`tD�\����0���q盥CB/іi�jA��۽B&��	����v��Ki���_��d�-K�eɏd����1z���N?r�	���ЀY/=���+�#߲e�!>����Cz�V؆�~��� Aʡ@�2ޯ}�kvX�x��մX2I2��SO=-���7Map�8��֪R��$������T���=w��wOU$_��Wl<|s��+���j����a�ϮK��1���^���J�^Xb���c�� �z��9�Ƹbň��%K�!l�.�BT���}�[�Q<��n��Ds (憹g|x>�q�>�5ς렐�ӝ;����X=��ɀ������A��D<s��W�#�M9�t	�%�PD4�Q�e={�י[��(�R��#�� y�~�:����,�����1<�q^gk9&_Y2e��7���g�c4�P��A��L�e�29l�(��w��(D{�B��nDH���E�|˸.пx�e`�ԚO��ڡU,{Wq.��;�E�d-X$���{x�\�9ܛ�Q���R����V��NcA��@�$a�7�`a��*z�x�y�Љ*��k��$� &�F3���Yw�K�da�p<^0DB>���,-��Ij�\#���A�,	y���UBY��&`�?����*���tSSr�M�w0'/���Z�S*�ge��	2��$�Ԭ�B9Wo����*���zz�dt�6ɥ����_6ޠ뮿Zb��F{�ԛV*�K}�fC�=�7���>+�C�<���w���f�Y;"V���[�x���3���uU������(�Ɗ'������f��Z�n��e�&찚����$A\��-�J2�H�ri]�0�1���9<<d�?}��D��B#䫑���gkd��j��!z8�n�����mI��y�!��`�=�	W�����`_���f�f �QF�N}o[��)<��,O�y� nP:�b%,�/��D)�رծ�X�c��ᢌ�ݪ�0����y�Ob��2�y���{d}}E�
�������U�V���L��J�~�����Ѻ�k,��9��)��;p�r۟^��B$`w���N����uM���I�����3(vE	�	�ڤ�W��VQL8�Ϣ0��	���Kw�8��ą)��s�-ܰ՝5�n�����PH�Z�q�jx��+�����Z��
ޗ���|�e��8-{vn���������1u�T��?7-'O��x*-1��z $�[�y�*b�˖c���{Ú��sֹ��J#Q�*œfE½RFD��8��_�d2�[n��/�ʙ��Ț�)پg�l�է���YY��O�-J�*�*7��}^ԈVwqHz�GժX4�K�⮜*�VcN�Z[FE����Z�Y�sMt쫸8-�ފ${f�[�2�;dIa*F�j�Y�5@!��A�R�����\}�U�w��j�?gm��th�:�Ww���ə���gܮav3�h!��PD��R�;,4'�*&��m�	��猑
G�9: Ⲭ�ͻ���W:*�Nd�;���	�+��R.J�y�T��ݻw�� ��*�:�;�;������H�!"�Q�8I����Ēdz�r�3�u���	U�!_�Dm 9!D�����	~^�C�X��fmP�x��E]܎������ղ�(2�����}E�CҸ�����y����=�{�N�=��3�_���?���l!r��y��߹g�V��R-�����n�ݥ/�}\ױ�kz��x2Ynw��!�WB?
c�,m��Vi:�y�箶pn��݃|X�Z����p�ؾ�#�c">&y�"���Ӂ���D�Q��-+�h�4$�
�Y+ꃕ�"7fT-�`kP`d^RSʴ Q�?�S��7�Ep��*Z�)%,y�,7����=O���P�X4O��t��ެ4����d��E�5���Z�9�� -� j�l��\�������P��a��旤8���dh�nNu5:AAV�0k>�ba�YzO�3�y��N�Q�v��F��4+y)�j�3�s��kk�H�Ї��X�B��� I�]_��r�~�Gv��e�O_M�c��������B�Q��+��D.aE�G��-��Px��8j��vۭz�V�"�O�%�!ްa�]o9S5�f�õ�B�c�}�Ta�	kLI;n�{��`�Y�qy����!f��#�z��������𾮊�g#L�[n2A��C�9��4z�X3����/��6V�l6R���H�ɩ	y��ˮ3����p� (VO����oA�{�����w�r�v.\�����}g(*��5o���1a�?���v-�
	��66�I�EM|oO�{�6F�e��nJ�n�_���~�u�F�Z����,Ð	Ϩ�X�^�O�[��[�r�"�^q�qk����44a�7��)��9���f���o�~��Qf��wU��<+�5��۲X,���R���Z��y�z�Ϫ���	p�H�f�,VP&����$QW&�<ua�wA,�K���.Ŝ�w:/l��U��iW��b���dp��Z"R�U��K'^��٠h�HJ��Z�YX,D���"�{b�f�(����h�I��sl(��| Y�Vp�h�x�k�ARy�$:G�w��I��7m�֠�T7��T:f�@K��S�*r��<I����JժKA-�Hݳg��=�ρ��W�b,Y�tA�~�j+BP3��n���+W�Z�,�}���M �n~��������F|6>�������_N�8.7�7����@]Lׇ�<!X Kk2��̝w���"
g8K�h��v��c,�>��|�_2$�>X�|qͥ��C�q�`�#x�= L����/h"�n�o*�''�\�Y-I�r�b�m��X�A1w��a�ؼ6C�tw�C^�����W��=�ʳPB��CH��]u��j[w�Y�����;��G���p���0��t\�������T����r}~8��WDgb�,�Y��x.����b�֬����J�e��7�Q~<ڧu� �Č��+�`�Y�B/n�3)���eZ�Q#�(�/���}8 y��N��Z�9�#B��ʢFg��c\�K�yч��
�QPj�-ʖX&��bN�ӼZ�NӺE&��ju��)fa_J��(r��*w���k�����d��o�]Z�
+�x��W�Ro��L��T�e��7k�	t}��R��GK�P�tL�7J�ɥd�ӫ֤^xV��U�����Z޼dS˻pn�@	*	6��"�b�*��ΰ*	[1zܸo�\*�X1���W\.�*���կ��?h��7�tH���Iss��������}jaΆ��Ç��F�`y�pTc�FH�>�}�b�"9�w�5��'}l��L�gŊa[�8J��+�ո%>�咭�Ν�/���1�>\����{L(s�8˞k3��d�N�=����{nG����R�:la�����
���{�;�i����e�����Jo_���v�������<=ۘ�^�dL�l�~޷����9x�Jˉ�pF���S,;�ߌ�ݡ_8����w���n��	�< ��x�ۇ�<��Ͻ��-�g����7T�#�	�O'���pM����o��sj�����^����&�=��#��ޏ�P�cG�H�<-�	�p��\Y���m{9�|�N�u���� U>��7c풤�.�%֦-�+��xܠY�-'��Gi�񨋽1��FD<�(��|��ͅ�"���t���)�kD�
���q:��^��Ķ�z騜?}\Z����ƕ�@�Z��"}B��Md�I��k��>3�t��0l>�3���A�&&�_mG�@��C�{ح�l;��k��<�CK�}6�����PœPTt��>��е�ˏIr`X�-���G `[(�d��Co�N��I4���?#��dH-���A�2�j�4j��Rk��0-��Òɖ�vc�s	�K�%C�2��Z2��,[$��4B3S�UH�Pvք��F��Y�\�J	�<�����%�g8����3���q�<�<�Kx������͊�r%$���ulnCw�+�7@7�jOօk��#�zt�����ߚ7�k���0$S�.b����B��_��7,!�r���|
�|ӛ�hBf|ո)*��T/��D��³q@L@����3f�MBFP.�]�ڒzx8 ��>��f�#�V9�'��=�%{��cb>�$^y��]�%��A�����w�b}=ʦ�B�g�c�����==��C��[�y����Yh$�?.`��w�O��g��~�ʿ�z���Z(��yR;<'��s�Ψ����y~E���3�bi�y""��u\Wm�;�"ﺕ�7,@���y}��g?�����u(�n||����j�YT��0��q��p1�c��/i�8� &f}я̝h�:1�L���B. /�a����I�9MS��o��r�h�G�@�Ye�>��y�Q�&��j�j�Q)J;�:	�@�]�E�r������|s� ��fյ��ROH�E'FGun�H���0y�}#�����vg���xo	"̿�a��%zۖ E�@gڱ{�~L-��*�)�/��l�ȁ�[d���r����
+$a�Ð�Q����TOAG?!�C7��}WmݓR���$
k��\��C���Z9S�h�]������ӱ$�A����������|Q:��������_���e���'��h�����`���=l~���ݿ�2�|P��~��&$1>�����&�HR"�� (CxZ�Z����'��y�Ⱦ�(�nx�)�v��I�U�H	�|�@GA %�o=|4l)�d	c^7�t�����x�O|��4eE(����B⚗_~�Z�Wɽ��+����ۘ�ʙGPT�����Ԓ*�5V�066��*��~nư�<ǪUc����g�yڬ�[o�%"o���?.�Wek����ݺ5��'ׁ"��`��
��fQ4YnǸl�.'6=��C���ֻO�������j]*�/�����u�r^ Bߌ���}��ȇܬ�O؉mǎ�v�Ϝ���'�"���dd\����H�΁W(vf��y��G"�p��)l��������z�%���U*]����׭w� �Z�A@R��r�ɗ6���>��Q`�Ȧ<t� �j�V��� ��2�4��"ŖQ;
~Kjv����̲6�7�Źn_<	*r��2=qD֍�˺��b����Gb�O5�X�$R�K�dpt�(fTs[�G���j��H�n�.�fAՐ)o:����rs��H�fKAˇ�¢2�����[��)'��im�XX�몁c�H��+��!�̙#��+k�r����m;�g�*Ͽ$����)��v�Z�3�o=./>'2�"�a�ͩN='[��G�iZ�1}v3���T$�T�B��X"��_G�"G%EVR��E.:}e��ݭ����V��	y^��[�r�-P�\���>Ò�3�1��E�5�" ����,�tBX�x$v��o۶٬|(ʄ���!��pm/�S�B<�5� i[h�ԩ�V�x�؉���00��싡 f�e����)Ǎ6�*Ɨ�`�{pp@��]R�9���{<aG���<���M�E�1�(���Ӭv>���Y�o�,�͜����{y�����⺿�ۿm��w�" q�6 ��S����̔�!�P�gݟ��.Z^�{*cϨ�m�{pB$O��� �x}������#p����ܣ |�_^��Ni�ӄ��0@@�<��1�w�#�I,|Ƌ�þ�q�Kf3>�e˟�A�7�&����_a�Z�n�_K~��tldߞj%V./آۤА��p<��"�1�N�1|zۅ]��
6��>1_)�
���+r�n�!>�?h�@�3\QS7����c}R	��[�&W�E��@���U���4odq���u�KR-���u�3��Tj���������zKuc�T����ͨ���Ӫ'
����j��F<�E^J��D�XK�����f����yI���
;�6�X���1eE^՚�r�3o�1.W];%��1���	�����"�9���I.�3�g�u9{N��.�PK6�L[fΝ�5�v�mw$��X����8�%��1�X�E��m~���%}C�FG�K�٠x���&8��K��E�../I@�<�?7�|cx�\|!���7�5���������G@�>qe&Jea2�vH�ƃ"����:t�]��hZ'"����.���C�DB��R��b��0��zs�o���z�Cƍ3�^0�\t�Ch	w�q�_mMx�`�)�o�D/`��S�Oɞ=;�~���s�\�J\�V�9�Y%�WL�6m���^'�:yMNN��*��m�bIC��'O�ͪ0��K[�u�a/�4��:Jj����q����Ϯ���Ĵ������ޒ����<̱�����nʞ��J��|��iD�	3��F�n�ŋ��ϭp�x�d�}�������G젌�4�6�����)�;�E0V""<��sL(҅p.n�e���{�&YU��A���w_�?����4ͷN#D�[q	��Es-�H�9B�p��>y�~�I�	c� ��nꆶ��%I�nN�x�$L��R�%V?�NH��J�;��TL�0M�D�Z�;wXj�s�z�Z�jy�k-Pk��nmٲ�>;�g��ɚ��r�ʃ�ʱ��o>!`Q�mɤ陚��x۞���1��Y��G��o����<<���mڈ�/���|�Z�u���&���\C �0�A�����(2�=Q&˶���o;(�*rI��?#��&�f�@n�̤
��r���*W_3/�<��a� ��o����K27u��sS�uc�ˊ��Ei���2�
L���=���T8<� �)�H�������V����ܻkgx�U@	)��"F����U�L��&�d�c_�1g��p���ۛ3X�
^��ö�������ھ��_�5K����c��B�~���O���	-����@���<p��xND�Bo_��:0|Xs�����yw��N�7�6����=��Ck:����^?_������ė��cU\���oa�D�`g�7^<*�J���u=5�-8!�
Q'&'"�N�(��Ҋ)���e�l�=\��0���Ho}�7�/"�� *߶w�/5tc�,q�]nL4��}��wk���ɰA7{��=��*m�����O�}�{��M���Ri��!�E��y䜱�xi���k����K�l��Ї�(��}j$e����+j5�OL�k�Yٱs{�Xy�s����9���r��ҕMs�Z���q���$���-	�&��'l��0���v�&n�k��zSB��*���R+��s�^PAY���A�U:f�FoOB��y�hP ��{�����y��S1�X�V-K��a���$Ez�E��j@�1�-Ӷv"�g~]����B2�i�a|�&�}˼�?����[�D�<����)�9���˓(��EB����K>���yY��u�j��JlA���l}k��m�:�,���˫PI�2l�3�9��>�m����XfD�J�_$��
�i�
Lŉׯ����g��\�&5P�w�]8�Urr�H�v^��;3�	lݖ%^�x�5v��f$������a��>s�����amY�Ř,{l<X�޺����J�{Vul��.��ܸ�������X�hU�VM(ћ*[�e�X2��c�t>�'�b�h�
��@�8Z���*b�L�9B�J�+��E�3���x��=V��y�K�=�R�1�X�G��b#�l��@Q�߹���|�ye>}�_����pl��"w��m�.����0/��9B���.`�kܞ�G�(c'��Ц��l����];�K�^M,�d|x���弡F$$�y��k�4��K^����U~��k �ja�Z�Jl�܄lۼE�U�ܕEhM�.	��j�E�v!B�JZ_�&J�1�^�	��]�G���S��Z��t²����p8��C���c�A*�i�*�v3t�H�&]����� L3#��)L�g����zГp��+�lK�`��-,޾L���iq���
��
�2���d�k0��!�ߨ�a�.�C�p�M��"��y(�0��F�����nU���P�κQ�����
{<)�Qn4C�Z*����\�U+U����q`�ɬ
�TV:FLVTA�`�(h��3�������Q�ɔ��K�N+�sָ�{`��ᵩX����
�a�Pʕ��
֍M����Ī6�8$Bkt�!X#���������~V��'�:��?/xx^�.G�P�� 4��r,�;wn��]��`���"�W�Xe��Xp�٥����Ș�y;�<|���RTے v�z�N*lW��ph,����ӊ��ykDO��Ӌ���:V��$�w����G�A�-�*�V��|�du0�Ldy�B!��u\�۞#VO�����`��?���PΌ��_:)�<Z���~̙�)0G$�}g*�@�8x
�	{<#BF>��?�㗽�n�{�������ɛ�5eW��pF {<��;�/��=�St4��x�o��z�}���q��޾(a��DZ���֙�d�yd��XN�rwf�Lk�'|]*�;�\��,'Z�W
%)-���5�Qf�S�>�����$�Wn�E�FK�x�(�Dے����
�GU��l�EI%;*d�j��%���)�2�z]b�j*�j��f)��[���SW��$=9�ډ�/���kL�%�(��i�}�\��쳝DI*z�x�c�(&��wH��n�Y�a��+r~zR�`�ʘQ�Zh��~���v��u>"zԴ��q��eIZ��I�tͮA�c�:���M���q��]o��
�]�K�f�ŲYw�%=x}���F��7�di!.�%�k�׭>S��,�	����?l�m_iS�24�J��+g^����ʉS�r��$��z׻���xFZz��%��K���Z),��_rVu2k��Qr1�%U��ɦ�����ܢ
's�u^zҹ��s��T����zK��$���u05-B�[�N)�x�x�K�xuBzݖyDr�"$��uW�"�?x����C���G0��B�_bڜ��^x�`�<xy��_�
e�X�+f-�SDC���e���g����bU� �������?&�?���q�ilݶ��X�	����cG�\u�
{&��r�5Ξ9+_��W�kضu��:6��}�I�>tr�u׫E�6}&�<����d�~�P��ʖ�ۥo�_�dvnV�z�iK��Gٻ{�QC3v��P�X��?��]oϞ}�CEb�/:��~���8��e��sG�{��2���R��ʎ��� �D: ��oz����?��O����}p�L��"����������h��T2eg#ފ`�bXLc�$��������0[�D��~��5�~|Ug�|�F��T(Ja��L�~EV��ȶ�u@��g���^L-d5��so�`v�DJ�qf7e��9J(Y(}��Nf��Ú�K�⛾�*1ղ\�W�X{�XC-U�歲4Ku���iwx,��4�KPd����͞V�tR&ϼ$��,��j���+�/Z�T�q�U������U��?V���BM\�C���&��%�NEdht0��Q��Uᴸ����a�c�q	{��S����^n��1��j��b�t6�j����a��<-F�	�6e]�δ �uT�C���y��#�U���������V��eW�G�.K>�
��UK�.u�3��L���l[NAn�
z�����\�c�>y�(��̯HV����c3n��&�Ԇ4�Q��M�\��r�Y,6�0�p	��㦩F]��UԈ����	)�J��'>�	;\T�(\'�I���M "���o�a%�I/Wx�;-ǣ����&���Iv2,�_��_�k��R.LLYb��`�r/
�I������8�����70�g�$]s���Q��2�/ ]��9�}�q��X����944l��T��_3��5P��9�H�.�{߻׼<��-�ܢ�y�]��
�z�����'<��q� A�o����O�5�W�ڰyX9>j��{�}?�g&����,�DR�Șx�������&Kp�����@j�|Z�%��{�ʿ$��Q�c��(C�n�W�v相9�9<�+��/�|@>��?���{Dab��v��
���6Ç]����X}��ES��O4w.
�t'^C:���y��M�A<VZ\4�$@��9��^��}������J�c26>(5+��Xk��=4�7
�͘TM�]�"�fe@]�lzX����5Ǎae�h)>Z(D0�K�ଛ���x|�b�踖����9�4*�jɞ��Wd�B �O�SK_�����h��{��l���#|3��C��n&(�V=��Ì�֗�$.�ŢJ�3t/Rо(�Z��a��tqx��iHO6i���X'�tb��Ĵ���Kq�-�?<!O?U�ӧ���==3�o��`5�i���M���\=�&})6�zoy�����b-�DhR���t+��q��3祩k���^�Ƞ���@L��R�֣~��8� �'B&?&�&�%���W�s%�
���n�s�v�=ݰ1=���3P t:����@
t�/���j��C��*}2�U���p�i]���,a82<f]�H��ܯ��ʕ�"b֤���Rܬh�^�Ů���k�戧BpB������[`���{�ѐq�=�l�*�e �
k}�U�˪��
�E��(����Z��[����y׻l>A'��k�B���R{��[�� кf\"��#!����;��s۶�*��ٽ���Cj��p	q�y��)g�C7�~�Ö�V�8T��IN��=x$5�a�z�Cx.���\����CɂB�2^��E�[(�gP-��t,��|�O�Ԟ���ɟ�{J�Οz�'�����ı\F9�n�iX���/���Q~��F���a����$^f�F�ϥU��Ӵ�׳�Ey�U��)`dy�:�=	ٴc����ftST��T0����ɐTKI���Tǻ]S�;�eÖ�r~�5�f�" p�\�����K�^�,����� ��n5�n���3Ν:�ߧdͪa���w���!��J�TS��>�{��,'�h�
�j~�O�%E@Z�����꤁�%[��Ե���n��Ta\��Nw5�k_fMX��Kx��'E�Ӳ���|E�J�&�r��Y�qD�׍KY-#i리�a<2!�^�j���5�BiVN�(����u{N�cK�j�Jdm���X!���*�<����'����������N����q��65ֲ#�jY���Z���M���ጅ���[��s�x+��`��{r=*������lK�k����U@�,|�+A�B��X�ZV���=�raa����>a�ݻwX8��ǟ	�I��+64ѴH�%������L�t�G|�Kl<��L�O�>O���5��G�Y'�Q
��o��F"=A����,�Z����v���z��5�.UM�?��r�=��},�B9bgd�����.���t_M������]��<7�x(sG��̇dr��3X��a=��[l]��L�aM�l��ŋ2F����衹��c�G�P��������2�(^�궐c���Ds�!�|Q�}Ȟ�;m�%�:�e·�^�/���<�u�r�/�it��|��������)��5�;��ƤV.JF7݄��U�N�<lŪ�c&��5�MA�n�@_BrJ*)cG��a��LL&�/��ܖLP�D�**$�rX�*��*�ә�Z�C��gsCҕ��]Ө���j,��|A�&�[�d07���WZ�����3�-(:�����Mx:�>A�cá(�Z���:X����Ú��%c<4��f!&�Z?ڊ�h�&�,#��7��vq��H�����j9��a���v��5�r��N���_���C$rÍ�r��oVA�����S���Ge��}VG��2Y��!#��(�:O	U�=:���K2�����������.�׿~�|ﾣ�T�r`t��E���
T�l-J�yA�I�B�D=
�ؼt��@�A��w�ۄ�g?�����w�-j��-1�0L8�i�X�ɉ��Z��=��9s���/�By�aٹ�5f�
]���;n��B	l����ǎ�UW�7K��=��J�n�:J¢wϞ��q=��}V��
%���808lm#}�;I[��9��|���U��$��D�sF����������(�]�vژ|3:8�[�B�̽�z�*=;Iko����"eE{��V��b#P�������#h#�͵]��э��e�e�\�ZŚǠ0�����D1_�ݫ&���<�ؙ�>77o�����a�,�|!�������P���o1;X取}̱�H�����^�m%�]4�V��G�7&U��G}�jx�>��?�#������1��׮��<uCX-��^�-������xE�)��4c��͒ǟR�xg�$j���&N�
��zǹBE�����?���
�^uMt�t'Ϋ�V!���]f�,�=_%np��*��^�=9�p��Z��,Fގ놯�PAM[>
g`(2>��UZF�c��2؟��|�n�pU ����'m�5����840l�Hx�x67T�Ȉ8\�t�5�.U۲PRwQ��NS
����rN�[��eq\�	Q���ݡ���%�]�!�q�>����ѓ�^��G��~�V�����I�$�2:�U!3��K�q�.�ˮ�$�k����A�z������,�"�N8j��Ւ�,����U7l�4Cņ��ڪ����\�U�����A�/�Dp8�w+�R���\��DTq� �D�`ac�:DD��u5V�����	����%и7���Dp�	Sҹ�,Y��{aq--5T�=1V"��w�U�w鱆9�!"z�u�u�vyA���)�V��"x9#,o�ٍkǊ��2.���Oı]���	��l7w�tV"�h��u��B0��T��V��`�0a��䱜i
ΚA�@���L���K�D�����[�u�?n^�j~O�ݯ�֛O�̬C�𳇹�C��g�`����R����ό��!��|z�f���Q/���{�^������⁺D}=Ln'M�P���s�U�4,���;VS���e"_�8�5��=[O�WP��_�ٸ���������$�s��]S+%Hv�m ;���z�Y��Lf�B�# |f�5UC�RA[T����,��s?��3��f��
Qbzp�e�����W˦QkOy;ޖ�
�x�rE-����}�x^6�����wmS<5�t0N����y���;@��u���U����3P�t"0$P��K�)��[�д[X����_΂ ��8�e�m�1�I~c�����t:!wM˰�&���m�eі\~��A����V�#�7�IJ��̻~����j�@8�˻�,[hz���<��5����0���sԀ�&��6�PewN-��1��dh�W���[$�j���)�#���T;5)����� 8N�8)c#�,�ΆM�Up.��K�'�� lQ����!�M�STҖ͕Tx��LH�\�s=N4\��s����X��v��mW��5oO>iy��Yי��l�0�X����G���o}GΜ=/�KR\t[�'�T��FY��&��5�8hcH8e����������r�� tתr�b2�OpH��qQ��x�w��y��jh��%<���;����θ&����4���(���}�~y���L9'��=ց��t<�7n���!�k�UI�ꁌ��Z�fHv��Uc2�b�<)���44�� ��(�}21RP��c��۶� yا.$�=�;�x#�0�<eW]��^�蛰�_���ˑ��G�]%���[8�}¾"���֑x*�w�P��2\��:��U���t��_�Rٳ�OU����3��T��	*�뭋�U�Q*���E��z���Mo�W�өf���=gaI-y���F[���DÒ���kKU�*T.R���P?_}�4k*�s�]8hj��V�E�ã���j���b����S0���(�9�>IٰnH֬�K�_3A���  ��IDAT���;4��ҟW�����-A�r,�$-���+ȂZA�	�J�y)6p�s*�v��Ԏ�ID:Aٸy"�jǪP�#�^fٓe�]dY#;����3l�`}j; $@ۿ�#�x2ĠGZM��-PtN���H�%��Kv8
�9��8�K������{D����Po%	�� ]m���NZ�J�(�L�BU��S%y�*���s�\7s�!b�����.:�֌=�8�]�}}�iB�?�O(1W.�g�� B�z�>^�+����ͽ�>���x1���E����k}���"�1ca�����q�J���t=��/=F��Ŭj�>��<���q"䙛��Y��������f���t�V-��#G|��Ysm�"A��v�m!�V,B\9�a֦G�0_F���ªt)�h^���g�PO?����B�>���Qr����(`U�D��'���ƃ������I���,t����Ady1&��#/�d�ֈ}Q�9���EI���OX/{�m�qּ�oG��W��g�[���QD̏��xO��w}�ӟ�����?V/�Z�r��.�o�y��IG���F:e�Ha]�,a�F�B,(�~��kb�V#ެW�mM:�i�|�k4�0����NCQ��Rj�+:NS� �9�M���p&ea��}M��^^�Ճ�͸N�*�O�X��т��{�o n�b�jfRMcx���Z�Kk~Rff-S����s	�c$��*-���%������ Ӕd�bc����jғq�'C�H�9Y�L��D��6s�o���s�\ƽ��≸a���B��z���X� B�s`�-4�`�޸�9� 4x�f;�T�y�<��q�y/�c>��R�Tx��r1�*�S�ud�Ԥ~aR�������1�~/A��;�]���%~�F�?�AJ'����r��Z\���7\��8/O�8)ǎ/H'��Ϳ{�^����G�x�� �h�Pr�ɸ)F���"��C=W/d|�?$^8gͺ�D�|+�A/�{�sp����6}^�h�01J�/��͡EQYBU�Kr����0�8dљH@�F�;����>{��Ql�Wl:��Bw�C/ y�v�T�|���(|��D(&;m+l�R9k�a��K��X��ѣ��o��oL#���7��~�<��kW�_��lH�Ւ-[6��6�u�d���'?��]w�)xGQ����ߓ�~�y��T	ߢc�5
c�Â��� �-�Qq<���`ɣh}��z��zy�s����uǵ�Ţ�/�T��sH>�]�V��B�������c:����\�®Ø\��֙=H��#���b08�<��N#�ĢC7�ǣ���׹M��>�5���6 �xB�\���T�`y# ���KVN��R��п�UK�Ԫ�2��VE�� 9�r���նTM���{�M\��Z���z�EU$�v�0�z����&dt�W�{B�H�j���W�ts���m�̝4��������(
Rx!I�jK;0W��B�7��Q�-9��R*�{2MI���m�]qO,��᠄�@�d�+zr����N����Z���	)\#��=�|G��j��޾a9u�<��a�pVdǮ�R\���ϟ�t�"�_�K2�Wsy�����oO� �|N߻#-{��Q�qR�mέA��*C��0��֓�J��[�d�¹��:I?Q�p�$���9��������Y�<Bko���&$|�B`�RkQ'%�@�|2�j��9ݖ���<!���{�,:P�ʯ��1)R`Cܝ1yk�ԩs�<��|���,v��:ss��t�� @��A� ��R��Cf7�C����uϞ]��$!����-�֭[k��y{�}�9�p��!U��=��Rzb�v�B�����$l#�^�����Z���˜���qVqL6oY��򮐒@�9�VH�� ăG!쮹�j�.��3j�
�r�ث���b&�چЇ�u FɿY�Ç_5e�Q������Ike����5JF
��}/��%�n-+�nb4gи��>VQ��5:���'�LB}�=��3�j帅��K��7���-cc��/�3!��F�ʵ�/�H]aߒ�C%�H�R�!�a��S)W2x�E�2�?��O�.�:0ς!��A)�L�˂���h���[Q�y�5�!���bR�vI-aո*h�Z���;L@ZJ��JFf�2��1*8�YZ����V��bt���n�R�%�&
r�dU�M�!F��K�z���!��
q1�e�c�jԚV����">\Ly�k��J�EΘ�-W0g�%�A��],���vܳ/'R.�t��_������1# L���5� ݈ɳ��_�̃NJb͔fE�uy��R�)�v�\����gV�).��qs��nPK��3��ϯ�1����e5'�?y^��͓��ݴe@��s�&���m�+[r�I)�VR�>��)��]{-���7`��Z��-�1�k_˅�<<��pa"��5�^i��kq����)��G�pQ2!��~E� ��z�K�;p6�3g�{��㈃�\9f(��_>,_����I`��Wȵ�^m���gBx�.K�(�{�@�%V�0}�5ay�Bb\��5��f��h&��~��_�9���~���������G�̰ƽ���<F?�J��NSX���9rԔ�c���r�3�/~�
���u����I�c�v�ω�i��\���]�wD��+�ւ����Xn��A�����?`
�=�~����'�}�s᭐��>�=��[�-z��<��2�|w����'���ܞ�;��̥0�2��X�|��(9���q���k��cqq���C}Cz`SZ\�%y��l���d���lwױn!�w]��Ҋu��W�R3��Kg(V�Uw��P˴t0UtK���-�߲���f=	uI*U#�ʨ��aȆ�֜%Iآ�[D�N]|*Dc�������eQX�с���$L�������Sy�ؒz	"�֩V�t��Q�&��<�F[����>HHa^M[�I*���/Z��]�!�R���Eِ�}_Z��FՒ�����ڢ�)H����}�ZIќ��)�#��6�߄>�z����k��̍�i��:��c��}�>�ˢV�㶇�n=H)[1�z�r9���<�W���L��{�j�?$����%@ t�A$)�<գ������K���dfZd�z�W\�M�;���$?�ڬ��_yF*�y��w�
���}��י u̍��u��eE�qjB��$n��s�`U���(>���%���n�,�������os���#���$y�<=�'���G�8���ƻnzq��)�r�m�31Z��V�B�W����ksĢ}���*m�Ɖ��UG�8ָ~��>��s���$��yn�A�0\((�~�ԝ<Ċ�+��WM̘y��	�8�N�Ӥ|�;���zE���cW<v܅:�{�c�Xha�M�@E�s�ڵM&.LXr�/y�^r�#Bܣ�4MY�n�)^B���̼1�9��>g����w��{��\�>t�9��$�&�h�.���W���_-����)����m|xKTOo�������'���S<�X�BC~�b���X�"�����X�q�<?&���Y�g�K��|q�Z�)�fm����0�ik7Q QJ��a��,��4:� �,�4�5|&�v��DNfqቊ
T,�>銢���Ɏmkm���,�8}vAf
"�~R�i�!J�/ʂV}�*�{{��Ҩ�	��BAW-&����T�i��N�� H"C^֎�-���2?��O-�\_�
�0�j,"�Z�1i��a=ƥnWWDd=8�Rw�C���*{��4)�\�I*��Ϗɵo�%+V�٧&�������ʝr��ۥR8+U=ă��[�+�=r��Z��vvo���TA�UC�)�)ݣOY7k=N�)ٱ�)�vϾu�?W%~A���"=����&$;z@v]q���È@ھs��"R�V��w@$�X�o�k�ټ���E65�@�0X{�IG;$�r�x,NG��ca�B�l��z3++�W����U`����#��,O<��LL^���\m�ԅiY�j�UyBmL\�s�k�=(k֎q���yP�Q���=�.�c��P={����Li!`��J�}�=����gesn��6s��	�v�� �',��y��wGmՀ��"@]�a
�D&�H7S#��?��?1~���E�;a�x�_���/�?��?�����_u����B#t������n̩����LM�ȑï���{�t����鳦�����[��6ٲe�y`��<���K��1�����J���!KO~���F{w
��?ʉ�p��o� �}�������B?��޽]�õ�^���s�����==޿V�EByIt���ʿ|�K�Yo$�5J�_�pM���:�O����һe��U��=�5����&lbj^ʋ�DϤ��u��Yt΄�ba��̻�X@"���M՝A�T�nL%�\�}�*�wM*��gK23W����޿^n���<#=_��:4L_Vg�W.L�b%z��Mݤ���ԭ*��hY��hw
�\9���ޜ.�n��Z��i����Q�LKE��T���˪�	�w�7!$#&J6v+lG�4|��B�����%�#Zo���Z�
ޘu�r����)UF�s�u�4d�ꕲa�N)t�EY�~X�.�,��X�}#֪.
�$єW��Ǎ6�|�yS�R�u�p��*�2�]��,�wsaR,����2��Ҝ�]�]\>"��8g���%���w�Knx�!��p@}�36;�X$���p���ja[��^w\��,T(#xy���ɟ���=|H���P��+�$�L�� b�|��!6V�;���Z�s300��l�
e߾�&�jA���6�3��3�������Z~�3�[�I��<?�x�f�d�=�#)I!T"�B��Gb����	P愊W�x�ծ_��,�V��yp{�A
G=�����a�@���$���[��OP4���7�# �DB�/��V�7~�7LY9��㎷Y����IC���x�)d���w����1�YA R1���Z�,qo�7(�n+�CO��"�Kä�w��O/��E�3��#��X=l��NN�>i�9>;���}��ya/���qox��}� �O���I�{6�m��ȳ��5�I�ʵJ��zw?����	�f�˥���r_2�W�8�-Ua��	y���\ap�Z�t��O�t��tV-�1��f^i��X�Lr2mq�B�B D'$&�Xt�2:���U���PlX�Κ6����j� �$[I��mK�`��V^N���W��P_ڒ'E���p�d�T�X����� oz���U�(=z��i�m�m-�VK��T�5�q'^F��E�]���Ktn�'\�\ё.|���Ęk��A��<P�7�??��3���G�[yc|�>W����t��)�:ߔk��V6_�^.��|衧��O=��A�l��" ��ڭ�ϒ�W�W6�����܀l�ާjQ�V��K��^�E�7#�w��gN<c1�u��E�[���$SN`�t�s��=P<'�s�ᣏ|�#&���O��~���[o�C�E�Ah/+�v�T����	�������g,,o������8�P���� �5|��Xaf��-r��{U��.��e3�'��я~T��A=�I�7[�Tgu�LXp_��nG�^��2_�wlF�4����>�;v<�1���9PJ$SN\aν��J a��P�c��g\1!5x��S,�}I�ҥ��Ay�7�7����෡�3W�l�_�oߡ�{��?�տc�������e�0u_oV�i�̖`�|�aS�N�L	go���
`�x�#�2s(�Z�;�#a��i��2���^U&�kq{�㵐����.,y���yz���m1(����X�G
�Vut��/���P]��Fȶ��p����Ԭ������@�ު��UB>�h�r%]����Yi.��7w��V�5�p!��
{tЇ�Q�֧£m|��MJ�3�2>;ɸ
�@-�R]2=q�E���F����Y��e�Ϟ=����4îm���
H��*���5���4^��)	!Rj�KR��!��|B�'m��A���3R*/I")��!��қ�I��	rդ�Ob�X�VL��X:^X�C�XK?+rjUA���ƜuuC1NB\�������o�N`W��g���F�Z��0^H\�u��Ͱ������9!ji�es1%�N���ce�oY.?�'�dƪ{�eڜ�%��WEMaYN-)�.�<�#�]����ڹ]�YhE+��J�)!�v쐃�Y����,��&]�
K�..�F bE:�iȄ:�����c�S���{�cb�&�C��U�:���z�������>X�(.���xP(`Q�r�m�}�fCUf����dR��!�I��p� �������L$4�,��u]�K���X��*!��?G(-�L�\(�k��p��x"(BaX� �H��ڵ�~�����(4<�����3�ޞ����b��f>Hx�0'�3k�E�u�� ���}�Л�t�U��A H������!,���뿶�3�|�H²
�B�._�-Z��y�����Ȟ={�?��_7
�Z8xXs����p�,1��B.8!��a.��X������9N��*ԼE��/..D�K��xQ1>3=+�{�ݖ������W"X)pg��m9�9���`ak�*������A�O�lo�{d���V���x���������L:�nֳ-�����C�*s� �.kф����F-&�j2ؓ��� �tusV����&��K����Z9��lݼMFm���29qV�z	zڲy��[lobrVN-��`ΚQԚ���7= 3S*��6���j0O�@������+cnI�O�%�L��Kz�uM�Mc�$gP����0a���p����VŐyR��di�՛�R�b��s�7�KE�	�3�qש��������u���~��@��j��"�#��A���([�]��xEv�э=k�-��F�:Я�ˡ���+/�����#����$�����cjBf6a�4��p�"�9!7��U�����V}�6<
��r�hE�l�U�B-��f��1�T�z0_��}�e���(��;�#6l��پo'��e3�yg�������Ϩ�����|�_5Aޫ
����7�p}�c�-v�j�B�%(���a��E�6 OM|��%��C��	�/���;�A,}B�/? ���f���?'�����/���ѣ���7ɕW�L6f��?��ϫe�F����a��W����9� Sr����Ǟ�����Y�X��g�{ڄ�/��/�^�am�5�EGP��G(J69 �σ�%n���Dm�	/z<�i�S�6%�e}�M7[�����/|ዶ_��G��e��{�L9�{z��C�r��1��EJr�+f�Y���	�o�T.�Я���A����D�6����p�I�8ȳ)Epp
���L�\��L;�}�m<'��,{�5<�����F��e�nq�a�kؗ�t"4<:� ɳ@��f��y�8~�)��{kK�����o�5kV�gLx
�NY.w��&4� �Ƕ51
�&,���7E1�;��*˵�O�y�H�oڽ�]>3}����c�WR��b�c6Ɏ��Vh*P۠N��t��xĵ)~_�¬���礨L�>t��!����F��g�(��.�Z�ux��J�����s��"�<�U'�,����ҲztL��j���:�~97Q2���rY�RI�]�P��KZ�01�L}I�
H��� xT�}1�m����c)\�a�Q4b���k&��b3��S?mW%lny̗a;櫶oa�r�P���x�>0"06g�0)���7�V�r�����f��]7&�_� ���
~��F-��[7K��p��T�8̏>*�>"��N����q��k��@b5S�4to6{�/��&��R���BYV��ʪ�y��^��~ʄ'��R�rzC�j�$����;n���"�u�|s�y�w9\2�g���I=�\���9t\�������}���$y�}����^�5-�037+O>��}n��d֨e]"�ϑ�gԂ_�Z-��~���DE��F� ��X�$���t'F����9Y�'�(�>��0 L�{17���+�n��z�>���:,�.>���6/\�ꫯ4��^�F.aB��<3���:���u�-|��<#��k>>�RSN8�W�2F�W(,�"CA8p�=ק8��0vcŴf9�]�`>�$k`ء��xwO`w�)��'�y��m8���57/Z�-�M��w%͑dݱ}�%�׮]-?���,��ϘgD%,=��q �ZD� �*o|C�d��A�[���|Q�/��3�o�I�|g���X1�~�Т.@���a9�4iբ�A[ΊOdH��f�W�����â���d���(��ԄZnu�jm�Tj4j��{�j���#�v���e|�
ٺCǆaY�6���Oʫ�D�sD����)Gu�����\,j�-,�{�zd�4+z�SsR��1'��	v�Q��u�3�U�Я�{��-��1y���8���5F'�	-�dZ'�ԱD�+���+��	��o����2p&�;f�0�8��k�K5U��v|�ը������k��:G���4!_�0�.yU��xݒ��Y�N\�xIN��������q����OJn@=����0 k�/�ИX������5��UW���b�X�.���Dn��j��1��}z w�J�$�U1�3�X��r(l?�Ϋ����p�	%����!�1m!Â/-�UW^�uQI\���p.oH��o�G�-��[o�Ք �C�x�6l�dnzR}�+/�B�פ�Lx�":�hA�>�Ε���e/x�1B+��orA�����\�ȿQ�3�b��λ�vT��^�dT�M�]�
|<���<�A�6m4��k�W�PJ�\H_؅bB0{�������k��V�3���By��pC�,k8z@Ny�ʚ!�|e�ƍ�uN�Q���q�5������E��5_����u�o"��������ܔ�	Z�����2��ޣ�m�Z��7�3Z���IUzmK�ǀ`~�;߱�:��3���2��W�:������w��k����?��l��t���ᚉ�3�|�wGoo<KF���`.U̒�tR]�N�eM�u��\�2kP<�'�hZuG
��a�{�3�+v�T������������7J~8/��ML�Wϋ�ғ�Ez�\?��Z3!��b����s�֌����&e�����!X!�R=$۶l�5*< 횙��� �/{��dGz�	�̼y�-�Q(x�0�v�ې٤F�zhV�hB�ݘ��F�g�̗�_�	�VÑ��Њ�(��4�Ѝ�/_(�z��{���{뢺�C��LFTp�޼i�|�{�s�v�P�l�;ɫ)� W��d�,���k�P�Nj�e<} ����v�:)�����6���ql$\x�:�����6j�*�82������Յ�ZG�S9��ž�;(���F��RO_��q�f�����={����h�"�ۖ
���׊l$0��g]4�c�V�s�X����͖L�������(r|_Gڜvl��<�n)W�~U?��Í�u�G��"�=�� nX�����71&�,P >w��Iɕ��+���ǺT�h��;�愰U`F��.-.����=�	ڿwo�3�k2�Ӷ%��$~��3����G�r�(�y��=��h#z����uM�����㽺�*Q��HKi �Y'#�f��}k���՜��!���$�r00�L�iq7���{��·�t1Q����q�4��SO�W�k�ݽ*\�z��&	�5��倭�L/<������6�f�p+�k��~�C(����xX�@�E!^G]�i�d!.I�k,�0Ő!z}��ʾ���C�%���q��8}M�~�����j�::��ǁ����k�R����b0�bQiC��ՐE����@;m�Pj��dR+�_ܪKus_!:ق4�h�C1EB�xoJ��5��3�Gk�Z�eia)��b�#E�f+̒��������Q�{��U�J=G�k����J��j�xa�Ɇ�U���>>�6U��b\T3L�pI]9x��ږh��;��Wޡ�!41.�-�f�o�����@������}G�����/�:�0�¢�	�$����<'���pH�Q��>E�C�X��]SrD(��7�%*ڳo�*��x#_�Bn��Xu(C���<�._ÜHv�~>γ�ndC��i`(t���^�V�"bh�`v��-�����{j^�Y�<���0У����>����v^�AM�#~oFS���iыY[i˲jI܍�b��__W�Q�7�	 ��� u$*�$��DT�s$�G���JQ�LO� ���'ֽ���f����W�s������j ���8'm���퀋�s�ce�
?� O�T�A�Q�=E�K��\S%�h��4���'��S3��Z��H��e0FZS��ڑJ[��RR�㵍�5�s�L|'~���4K�]�V�?�:������k0՟��͙U��Q/�W������������ٻww�e�#�����#Bթm�dm�����k�m^���ǯp��>F�X��@��k�y;��K�D�-�M]��;�ź�x�@��BI���~�J#{�s�(]���p�G�(���1�&�b��5iԉDc��U+y��l�N>x/����ϽG~�g�T�R<�̖��>K�OO�6��pGc)Zgk	c�0b0�� 8�W��)�h�N8Æ̧]Z-1�A�Ԁ��բC�C���S)���)�8e�Q��x0�T�~!EF����,�m�m��R����"ܑ�sS�_��E�24�Ґ��BQ�PSl��ԄT/��B��Ϲ.Q��p�,W��k��Z�	�#T��b||!�`��؀�(��G%�xe�w��H_�+��{`���)�J�ׁ�CwS=$a��r��Bmj[�V��͡��v��Ů&��ñ-����FخYx��@��BP�Ւ�x�# �_V��i`О��h��߿$]�j4_P5��Z��q�Tm3\�,l�*Z���v�/�HiA5�k�wk��N��Ԕ�b�-����Ԯ�:4z�^�����n��<�=W�S�$l�������A�q�4$��yb��~���5ۆE��M�4���}:�����G���4m;}���c�^�fjiƉ�<����w�~�L�����(F��~j�ז�3	�8"'�z�n�µSirrQ�)�[p��)����qc]�b��R�l�5o��4��> ��^iC¯�|����r=O��P�\�;��=ԛ��k����6?C�=
�)	e@�,�#oL���Tԅ;�a-d�1�,M�BC䕏;,��/��3�/Qj��=�t��� .�H�Pa�\�	�:�K̙Mf��%�وX�q���4�Z&;:��^����@��� W��b�Uyi�(���������9WT�W��uE�C����νʸ[bZ��m)�]����NӐY��!�<�8k��LÔ(S��L?um�t�81�&2|�4�YV��ݛ��l�k�1Td�&����u��l��3�RMFq����#Vt+z2��B997*��DM�49��E��*�1D$d�b%��1p�X[��$�W���4�p�R�^ X.'�G��p���
y�RC��3g�	�cb��wE"蘃e�F	�y��C�Ǎ4�<�����e���C������cokT��8�W~�ȆnW�d�9<y_6�`Y�/��Q��CoP$�v@A6�S�h�Ct�T��;-s�H���U�'� ދ���*L�Z�Iߑi�{�a� C���r��֠/��,8 �z�Ҟ]��s�{p~�����78�R^<�CR��b~x�'�
C��Z*1my�����|�KR<�F{�:&4�Ԝ�F��d]���
�4�:c��]�۱j�O�����Ms�Y�V��{\��7U�G��cl�d .^�D���O��� GWYvޣ.��?��X�XG:R�W/*�~��9ZP�Upd�^g�X_K��� ;H�v7흀�i{�r��vk�`x$I��5r�|���i.Y�.��L�ox��vHh_o����-a4 ��Z/Q��P1, �^�@x_�9�={b|a�X�Ao�u�^~m�\��*_^��M0��<u.[g���-�H<�!��b��fVh��:����(a�+�����ʰ�k� � �5�T�X�$�M�RI7���G/֒�l�"�e����=1D�Wf���a|.���(�숾�몙�����hh����M?'�QF�y��۲i�Z��;3E�DQ�r�t�F��S��X2�0`�"�hP�:C����2ia���!�ru�~���iz�G���,��VX+���'�������~�R��(�k?UsE������iz��w���&���L��F����D�g�n@�`�t�����?��?�IPс��7�Fa�q8�����-z�G���������RCN�_����jEǫWg��Ek��aDW(�p w�R��dݸ�_S�A��w��Gj���
5�h���ik�Sw��C��;�[l��Ǳ7do�:mr�x ½UsEC�tK�7�S%x��<����qlڣ�޴�S����u�@�zOT��pܚ	��t$�9α��Wc��E��������D����>���;%|u4���fJO�\��@�������P�I�sϽ@����D�(#��|w�&�yxml;��k�l������x�z�����3���GNk>ʠ��2�1�tQ��rh�L���;M�}=Rp�W�|�вɳ��g�-��r�*���0;�٨�d��7��v�})�
���9z�i���|�`$R��z%�8���ش�ґʎ{��q�&�in*Go���X����&{���ea�1�O�S�1�\ h�����6��^VӮ8c��d�F�=K���vm}�=�4A*ك���ZM�:�VMQ(Q�	հ*]�0X������!?�<<_Ö�^БrLOB!�UW����������J�8G�kO�zG��x��J�iҲ$7���@�^X�*����g$�MK�sB�D�?n�k�r���ߛ8M]=K/���������� R�������x��؏9�F�$���C��O��<���U��~����O=D�L��O�����x��UBat�����;g��^`�Ǐ�
ݘ2*�r���I���Ģr����������2Ґ�w�{���=���I�F��)W�F�o�U����s���M?�Z������S�3��֟�i�]��@���P�8����<>���3�M���N��ǩ�&�*�l�w�hG�ht��h�_8��B�q�Y�Jhs�O;F�Chi�����nJ tn�ס�����z� ��+[�o u#Hj��7�-Q�
�"�66��5��S����ߥ�޴�=A @�i@ ;�N�i����s}?;�!���!�6Gʩ˗/�t[�%��\�n�����S�g������j��g�Q_�fT���º�@�4�m�ɚH1�ˌ˾�>zd|�?�#����A6���ݽ�2��Y�����ezS@dB�^��T� �+UOn2���-����@�$	0粘L�`a�T_ݠ��${�UIk�3&��)fv���T����	�|�m���h,,S��M56 nr���W@��F��8���e.��\����D�q���I�?��^�!�4HA���p����(���O���n��#o^��F �����F�)˨E\{t����1��	�8�z���'���d������ 7�J�F5��6F;w���C�|��;�b��l�5��%���^�ҵnC�����
�Ԉ � �U�4�������-M���Rd=w���A{�C��b`�'N�-��ꫯ����҃A����Dx��wx�������J#Ã�@�8��Q;�x�m�^��m��1�K�n��:��d��`�����و���+~n�%Hh��{����Y�;�&,tl_�x�	Y�p\�����q�Zь2ѫO�$]�T������J�l+T�Gj�k������L�nlÎ$�X�t*D+k�Ę'y�tc������$����I��7[A�*�o;і7�+m�&�R����ٳ��t��X���F�2�q��G	�|E�W-#� ��~S.|�Q���~>��-e���k"E]|\00��M���+W�d�V����<�g�,S�Vj|��&���C���|�:�� �*�`0�r(�B&�ˁ�{H����c�L���%���t+�~^LA̐m�� ��B�D�o�;c0	���>C^ϊ��XW�s��tQ���ձ�S�?E�����ߝ�=w��w�(��r�R J�{ظ��o�m	�2��P�ᐔ�0��|<�T�0�N�}��S������!^�W��ES�T��虗����<O�XF2<�h��������B;C�ylt�"����R��}�]��>�[x�R�p��ۙ�):pp�/��ea1����K�/о�{�8|��ߕ<{t���
��/ �L�B�@��o[�������u㌱e��sϧ����L>�`���n���t䤽z�*���o����R#���\�����$��gi��TA��ر#��9�s�~��N���O�v�{c��=X�����Nc��Q� ���M�0Gwή�U�Q��#�T����d��Y�ԓ���;A.4�A5-�KjT*4$���4��L+�qW����:�\��s�iz~��=��ׅ�UјA=6$���`/�׳��%����	|����;�vӁ�G(�^<�-���ڑ0��%�wb1n� �.w<�������u�,�&;�4lp),Fgǂ�b�2~^É {��Q�����i��z�^�
_)&��P�瀐�榨���e��pK�2�TZh�rD�9xW&�����ml�"\����%�V=�l��|=����eʕ|,&�w��P�])���e�UT;�����tN$쉏�;?|�����-�&�o*�(i ���_��)G��vb���!:s�gEwQ����UZXD�}�/tv�l��z�=�1�(�b#���U�O��A��uCM�æ)(�"�PVӁH�Д��CDx�d���j���9<,ccCt�|B8��S���������ݓ視"`��@���m�i۝���<�P�a�u=�
�0g4�"�������z�&�����A���}<��s�L��Z��c@�c�P~�$��i�����I�k�:N �����J�nc��C}}�咻��f���쩡��'�ۅ^��c!א4D~������^c�:$��B�E%<��c�k�.c˹��t��g��5��"���ein��MO
X-v�͠Gw�?D�8?��4���G���g�T���{�vV�͈@b!6 n�����AJ�q0�de-�Ƣ*s�q�A��|nX F�(b4)��t�b\a�C3� ��k$*� �biЌ�At�����}Ghf��2Aq	�p+�u����q&�aa��=�����4ћ���2G�To���h]ח��l.ӹ��l�uB
-�d�=�V�V�[t�j���Y�A�����6��it|GZ�R㈥Ҕ��R�cc��v ��P���}B�0�����T�++��76��0��ZC#���qz.*�+ ox�h��]$C�^��Ik�&����a����AV�p5"�<+�t1O7� oZ�V���w�'O��V�����~8ݎ��r��G4�Q��E��=?��ߚ���k��u GJ̟��ѳA:�&��D�/��<{�W�0�t$��l��Sc���e� 5��Q56]X���mI	v����U�� ��[���29cx�Z��l����X�vU`a��B%d'����0�2�Je�����4�W>�VM:H�����[Ϥ��Qi�G���8z���pG���RoBdI{��!\/�H7�{y�����W^~�����'v�Hg�L��dEI0�^g���	�>(��c��������\q���9p��!
ڒW�@�����,���[u>G� !`�LEyǿM' ��K}�$B8�ԋ) �E��tI	H#��l6�(�6H�ސO�Bz'ċ��`5;�HWٳ�J����*�ϭ�{﫮��W&id,C!6jA��CVTR[k����'h��N���� -@ҿ��K�ߏT��Aܬ��5�y����V��>�đ؆\WDf!BΑ���IG���!����?�F�h�Z�FK���������?�أ������̜�*�ȝkO^3(����!r������+�\2#'&�O{� p��a �#eT�)�9���죋���׆f&D
(�I3RP=���uہ��k��_N^��(3FH7Nu�=�W��屦z�a����422�`��;F��+���ǒ*��X�Zf�������9�1�X����3!J�����B�������<�>��@g<�d�h�R�6 $鹆59=+�8a�L�	Ј ���"��9�5�p�����
T�5bϨɞN3�h���t����.p��{xӡ8���NL~O�T���vu���E+IS��7Lt�����)������ a�<���	����@�F�����Hg8T�e�R�Sb $3^s�UbXx�J2���dD�m�����Cz�� _�[ڔ��(�"O�|��ˆx�������-��"�T��-��H�$zS�؈��jJ�i��.Հf��N���yZX z��t��$�e��:j��h��%�j�b�,���պO-r;Aޝ���E0r�� -�/���$�e������E�{*�
�!6ΡP����W�19��Z�NLI���� �8�LmL��So!?���h�C�K"����u��Z((�D�{���/��������������A�D���c��}5$#ަ��t�4ָj>������k�ap��Yۚ���?�v�9��kw3[���s�Y��{&�����z�y8M�z������*-/ϰя� �cǏҮ�459M�;Gym��}��$��W0 jh�J[��8?���TJu)k�%���'[m���Y���J���\�6�{��8�h"�\�S�]AL�lh����(]���xЁPPpo�sT�cJ��|�RsH���
I��q��g����((�%�a���(�v�s	�8%��'z�ѻib� ���/JT0~p� �aP��3��S�\���,R<iP�@ك5��B��'D��\lQ�����0{H,�W��d�n����Ste8	��.��*BmDϒ+3�tG��	C�i����&�oǘ?S�퉘�����m!1,�s_�L.�zg�#I�s��TZ��� ��'�2�BY��i���PYZ���)^�tב�t���
=��^�1���/�st�$l���"ǌ^�:�4�*+�1�1��911x5~H򅒜N���z]�j��ͣ?b~n�-�����Zw>"����"�@Zy�$Fb`�Gr��~*�x8�� ��=B�J�h��2�guuM*<�HA�r��g�C��
�att#m'4[��-hlz��i���|��k��nh���tCXXJ�l3��zB~c�C�O����[�<H�P�����S�g�Jx���IY+��z��Wd�]�t�����6����f�!�T��j��������x�:���wƮ	��@�)F��F0ؕ��
�Ikͩ2�5���5�v(�J��Y�5�i�l��<�k��+�A1�_�#-�`���iMjq�_ȳj���&�4y�HΨG�=D#�2tpO/-N����M&d>'����>���:��^��{b�5(lQ��c��ҥ3K���pâ�D�̥ͤSԕF[x��s��]��{z���irfI
�!4�T�mx�.E�����P)"��������ߪ�?����t��y��#N��	���J�`�*+M��5]��q���D�!����'2* _g���+���4���ӣRP���{.O���>��	a�	�g=t�俢��%ʮ48T��3Ν(6�-���R��%9b�{��P��N�j�a["���%M3��9B���-�H���3?�k�-iHC�fht���ۿC��2 㭷Έ$�"���ϋ�6ƪ���{W���w�(v����ӌ)P&E���#����)���QU�Ax�W:�]VUh�5(�(����;F�M�_�y�^b�7jn˖��=���ƙ�v{�̓�ߣ����mg���l��g+}ok����|�V#��;nm�7_����;ZbB�]���߾�g2�Bȶ{� �#Y�8�T2D׮�3�'h;�-��C�ig�2���5?�;JɸEk�e���9Z]^ɓ�m������O��l}��������un���6�M�G�{_�xM��ժ-n�t��I���T�1��>�󴁇���a`�bh�ϴ�]��'�&p��'�����V�c�y�|l���L�on�J��_{��F����?�dK{��l\�KSY�8k|A��*񃟡��_�4�"��I'�=�\�hy��`���kb�CԠ��5�l�֖V����([��/�AQ�J�v
�/Qݰ죣��JL��M<�}�ғ�����vOy����)wp��VW��K�P;�L�1�ugz(P�TG!�K>t�&v�
��Nʼ]\Ch���N!�6�=6�qP�V��^�Ɠ�� %�����S��sOP��[�ޒ\��`S\M���P4(�h^2@��f����w��Ō�u׮�B�*�8��|������WN����_��FB^x�����%Ճt͙3g}1<�����ȿ��2�-��������E�����NXԮ���D�M�d\X`ZdM�p$rs ��醭@t#`�
�������t����þ���c���a-��L�F%�1Lq:q�^A��g�/�����ٖ?�J,���uf�3�u�Jp80�����َ$:��:7�ߗ@0�P��y���i�|�Ҵ�`4`�%K�#�Ca�FT�����vxl�S!V�&M�\���*�I�:������``e�A��A��U�Ǧ ���JS<<O}�?��=�t��nz��R��b��j�0���n����:�O��P�Zf0/����[���7xo/߸�2�[tt�Q�	�!�Uq8e�U�ɟKC�K�:tlB���m85j��Ϋt@^$�=��Wk�������"~���񔖉'�_�uSJ��L��>0U
��a�s�GC4�c�QZ����z��Afwe9/L t�b���������w����?,�u�J�!�2���ʠ����9DM+%�@T�J�-,��DuLJ�7�&Rr�pV�^��:wO�]�Mz�hYg/�c�=�g�}�^y�U97��{{{�ͷ^]�/����-��7��U�!>u�B�<x�p��"��f�ve����C�b�ӟ��K��\+��ð@O^S�p���N5��Fi�[�%wz��1*n�w~�VAx��n=����a���E��>�5�;S5�AHG�����	��Y@:EGu������p+�-r��#�h��.Sʖ�������B���3u�M�5����u�#@���z�;���,���F�'jLċ,~�yq5��T-�%����Ɂ�i�lp��>zbEJo=��ń�u����t�֛��) Y��E�Ќ�E��Ñ^��O�E{�'hej�ν�@Fr����gD3���Q$��{ٰ��[%�7�@ZeeQW��οw��z}JB���ţ1in���lu����%����_��7�6�S"��8�	��d�g��j���n
 �6�͇J�QvR��&�����k�b$t<2�� �W�usLO�,���nd��o[��Q�7�q�dR���ư����I����� <�x"���D�XJ
E�c�T̑HM�4�;��!�V�Ƞ;8$�-��v�c������k�2�>x$����:~QQ��+�����A:��W��9>*���=uu���I��a P<m�U�B�ښ2x�@[�-��7r�Z#��9���*n�7%�Y�R�]x�è�l�u�(6��q��z�m�j���z��u�(C���d7�Zóǚ�&z5��2�#q��;R��dRRhWN�b<��ċg��0pN�ܫ��B[�"�t��\����Z^^g�J�f��˩���?�t�����cw�Bi��i[�RӐ����1dQ�MU@����%<�5B�+WZ�#�#��{~�� � �ԢJ�(����R��q�H��~�+�i���R�h�p�~�(����g��]#�����TO��������H���с=qJ�;>;}����<NW/��b�@��!�ޛ&v:���TW/-�l :ӕ�h���fg��wO0h8�~�P0QG�Z`�Tw��k��#=!���O�KX�VG(ftx���R8&��m�P dxmmypn�I,Ҧ��pʼP{/���=��� �gC8������P �KJ��Ý�{�)�D��W������7�����?8�ߓ��ɋ�X������%�!��H�	5��/ê��5QB��<sxC`��Ra��u�!���ڲ�J|��_���s2�L�s�ޣ�����f~a��?$7r��N�>#^׮�=��ÿ�
�T/��:*
�����D�#�$��߆>�D.��K�����t�V+ՌǎGŽ���	"[`��uz��}N�{l�ST�0l7��X��v���m7������a�nv�s c�Y�P�:#�g�w�w�瞕�qhh�VV &C���$�< ���%~#��t ��臔 
�]Mڊ
�R٘q���z�F���~j�^����SN��^��y�q����&z�A,��ժ0I�Ӧhh�#]R^\^��A��<Y���M�ӥ���)V2�-�#X9V $�9xU� @c�^]k��Gm�ʗ>K�J�~���e�ՕuJfثLb�K��L����Ը0�(�T�\�����I
g7{y^�l3D{vghf�q�;J�k+���ћ��҅��t�`��w�d2���mw���R0���
ޤh�X���j��ʕ���-�u�BD*��Ta�����b��$dH���\��G��K_y���w�Mg�Vh��GB�v��,dt[��|4�e�I��K�Fw����ôg�/��a;l<����Ѵ��Ű���㟣���N��d�X$##l`� ��w��)��ȗ#�ͤ�[u"�`�!�v 7�'���������~�=mt�NJ��'� !]����o���/K���Y���S`焂j��ǃ�A�N�>�S�@"O��� � ��ׇ�DEm�e��m+n؝�m����;I����57J?��v���������������s�z�R7(�+ o�""s}�'���E�v�S��Z�iA���jMQfE���C�֪�[��Ӄ�:�H��5��ܘo�![��ɀ��Y��M��U�b���<x�p*��e�@���Ү�8y*K�HE�bA
��mU4����œy�h���A_��,L��{�Iܻ�b�&-LM�����-�z���g�%�b�^hdV��	%��n��'�PoW@x�`��-~�	���E`Q_�`�-,�{�T�VT1�+:_���`U���ǖ�LA���J�up�geVwz�jn�k�_�z����	�)�@8"�ޓfC<w�H� ����������k�������Bi�A6-4���� �p0���1�d�酄iV��c�kR̊P�H�N=rT����*{݉���}�*4�k?��
����O�R�`��x�����2nq/{��>�������>���EJ��.��b���YwZ�@�~Ʌ7�F�:�^�����Å�\�a�F����~��P�WV����2T����u8??'ǉ��������3��$=�O�'-m>���὏��5�ܨ��|���������y^U�]x�z��i�m3n�FR.��5f<�7R|"���^�D�j}�6��zx	$=����q�b�Y�],���ג=�{����������G���:^'�G�w���r+�'y�Z⥧Su"`X�)��J�ܱ�����p��B!�u�#��m�mˣ*\^S�0d �z�*�
��ʖsi|$s��2�=>� <E���v��u[�X��^���@$K-7N./&N!� `M5L�^mI���软�im���?����C(��J�DH�MV�M���A�J�&��7E6��0)�ݘ5����&m2!�SIec����1��ǻ���t|=֧�a�ȵ�i�hye�±4�#�^�3t�2ѡ�=t�����X���&{�ْ���0�M��O�t��^]�W^��l����3�w�wd�ٓ�W_�B3�� ����-н��e<�a%e���;�ٗ)O��v6 &�.��_����o��z �F{ ��������K�O>B;'v\��P��1R>�L�YUQ��ӓP�@c�yz����ʀ�W^yY��Q��Sw���5�A�#�ڸ�B�m7Ƚ���	��u��N������b�/��|�Rϙ�c�����$�A��Ojil����A���55S3�P�c�p]N��vL���9��������~������A�2]3�k��²#2�\�2K���K�A��.:.�tA�'Ь�$O^����D �Xo���@����vI��}}�-W��P=��A��I�_�������A�$� &K�"1#{\6F�U<�sٛ��A���[�a�d�-� �����Zc�*|844�eQ������4ˀR�R��e�I(� ba|�!�(Q, Q��ᖩ�@$�B���q�-1����
�ޚ*�)v%f_چ)�� [���Iz�u��ر�k�5��>)��C�L�te!�b���U���x���
��a-����=o�NZ�������3*���5���2�Ok���� �M��F�V�k�7��>�����7e� ���	 W�|��L��a�Qؕ�_s<��?�^?�[�2ʈ�S)�<��!O��?��0�	k&�\BQ�'�����iKG1���}{%�.����o<X���~��u�(�?^rs�]U��z�L{���S�����>�עX�l
�a�az�N�i}�M���$=`D�O�wm5�9�N@l{����t�n_[S6[��F������>n�7�^}����5�QŦ�������Fӯ!֏����P� �l�K�A����]�fj� o�=�b��_�:��)~�2]��l䡪�hj���#��&�� �"%i,�y��s�L
���֢Z�!y-����޾��3Z��2;r�|�9����უt��Z���@S�	�B,��/5���m�]��-ѧ	a�_�a����A
Z�C�I�18495��*E�<[b��@��#]��4����l�󴼖��ǚ�	S���cmrt�s�����]���%3i}/L]!T 0fɶ�^���Fg�W/��!�F[kˡ��.:���:jQ<�S�sUgO� �fI�E<��ޞ��8u��b���)�����������9���چ�ך��w?x��'�Ѕ��t��ed��5�ƾ?�#��C��T��x�b|��¸�� ۳gA�U���� ����FaC<j��7���^9{PlQlŦ�����-a�`h8���F�=ws~~��k�H�\&�r���&�C�,��ޡPP��*����p:�����f%s�T?؏.��ȳ��U������?�s�q�Lz�9h~���60�iJz�R�v'�������Jڮ&�m���5r�޽��~��EZ[�K�ގe���x^��w[�M�5���J�So񁆰+��P�o6�Y�|�.4<՚��'�J�!���NZ�#FR$�'��.{�e�o�@UlK����ȽQ:q|7�,.�3?yQ�˻w�|.�[���'/��S����P5=i����'��7�����vN�1�� .��I��k�q���J�8��p����M��%��R�b����{F�R�8�7*�22�pERa%*��T8�fa*��S"�\���]_�5�#�B���t$rR�4$"(�������u�޿w�HW�E����X+
�%K����@��P��/t�.�Q2��k�@-3O��:�3!9�|n���w�X+M�.[���$,��b������$.�`ĐY��<����Q����l(>h���=U\/�Mn��� �O5Rc� �B�Ǆ���!�*���!:6j�rP�8��0n�f�\���Q�p�b���f;-�<��xmz���m>�M^_gק"L}Л��z(I����
���$3z٩�O��A�4��F�Vp�����g	����#t�c�
��nTSћz��{��gk����FQ�ֿu�y�@g��-l��-C&�����������[$��_������G���9�GZf�A�9~4K"!^́��vBi�	@���m���r����(L���M]� ��ǯӥMN���}�=���i�u��P{�I��]F�(�WU�t���A�t3���re�.^�a���xnPEN�����R"�%�P�a�<�G(��� ��	ZY/�B���a��C�E�NON%�MU|�C:��Tw��i�k���7�)ݴ�1�Y��2_�� �-��u�B,��q�VU8�r�������	r��ٲH	� �T�U}�c���Dp�\b�9�04�1W�����z@���>-���!��)y%���tk��9Y(<)m�--�R:���7�b���p(�B{.����@�����Vc�d0���{�)��J�k�;B�etg!>�}�n6е7咖@�`���a������iťߤ�m�4u�;RWz h�/>���QG���H�S���#��W�K~��Gg.�v'�������}���߶��7���x�k���k �C�/�������9t[�ٓ�v��L:�%S	~Ț���R�;<l�	�@{��n�_��Ҷ9�d�.���C����4�a���ㅬ�&����!����ߠ��4MO]���"m��~`� �.��ͷ����܅I:{fRr��=2j0	H>>d;�ޙ����&�y4]aqg�5i�ڵ/�߭�ݖ�Ρ+g)��ޞ�{WH�A��[�<|<� dn��BAr��қAj��P ��mB�"ס�t�C����<��(*��эrQ�n���x�<��9QC��RUr�����R�p�� �Q���DA�Q��l�
(��ɨ�q���L�b�#J�v�=�UW�P�')J���Qj�m
����g��	� �J�1D�B_��R�C��6ֳ�x}��*<^��P�oԶ���������;R9ȕ�Ԅ! O^ɔ�p�*�������jC�4���d{��ʍ�m� Y)U��ۺ��LU���c���z�U��y��B���;RYw�o}~���u@�;>���h�1��<ytK...HW��������Ll��0n�?�����7�[=�_��a��Q�;6������v�����{+��3]�����/
��<�6�'�s+e{y�h�u�W�kY�E)��	A����fW���&�0��
��`A�nND�`�\[�3Z�ٳ����:����_�;�e����[43���.��|����%iX�%-�҇\wO$�,gO���v�z3	a��,N��)Z�C�C��hhd���8�s�
����`�TB���KY���FV���Ӯ�(�WM���=@�wߧbݕ<4��_�Y~��b~�]B4K(�r�\A8L���B���|��	��Ď�'����4��2[ÈR��UV]�tq���"��?D��+C78����q��4ye��VJ��R[�=�F(JQ����T���Yt�ʴ���Z�� ��Ar����.��@S|/�����J���R���R�$��\~�̻lk��q��{tϽwӉ����~����N ������kY�F�7���K��SO�+<{�&~�7S�������֥�s~��yý{'�P������?���o�^
�x�>�D��|m\u�RK!Wٲ}��;�J����f
�E�����O���1y�G��m�A�AG��y��	�k v >i���g �h��t邀9@ǎGG)�赺�v�����0o�5@m��ں}���v@����s�x�u���ђ~kgZ�Է�v�F�Q��1}�����>ۺ��k�|<�pB�����5�Ih6-��:�)l<��%F�����&��ўLn�Wj��b`�vE$k��G)��}�3�Rw���4-_k��괼����R�����:����H4��7Ā�HA��mBͥb1G��]#Kv�&��PXl2(xu��҂�Ͱ�8�gP�f�f�����T�M����k�6��b�' CN�=Z��ؾ��p�q6��ϖ��st��ɻ�|%�`���H�D���8M�{����3T*�L�SO_�/}u�v��#צVh���5z�K47ET����Djj�v�즵�6�%J�Ҕ]-����i6�D_����� 뮑�=�6\���`C���UZ�K~��4=p��WT��b:�˯<O��ҁ�h��%�'�t������C��&<ӿ��Af�~�S�F�b+��B��6
����s��D�B^�Ј^x�E�A�^. �õkKB��q���g��^_K�C������u1T3��b���t��/0D�S�Qp` �^?/I�)Ӕt�V����@,IB��R0x�D ��;��?:$�:@� �?��0���,��w2i:���(U�y�?k���ܷ��n��3]�i��o-�vn��~;O��v�`}}=������o�f���sީ�d�m^�jR�0���^�󔜽O�-����^]f�Ry��V��:��E��T�hl̦O>v���=2�tjj�^~�-�Wœ��Y�89��c�L۠H8�@�R��%C@J(�Q�^�`�e^�A�[�Z���
�FzW��J�.졖�V���D�rC�` �`Ch�aɑBq[����[Wj�� ���[>^-�9�ގ!��s�tN�4Ǣ�\p��ӗ�=XH��xyIK6�ͻ�%�Ş:���Wk���if
:�+�q�V��eE��+��E)�e2���Š�F.I���
����қ���FSoY��KO�-O~��Nڽs�Fhiq��y�=� �tl��gd��i-�����Μ��:�4�b��c���h�u�/����^�3g�p�7& ��d(���T5�4;7-���!#mp������戃��%�a|ڤ�֐�SMi^�!��*�Ix�px`h0�3�Q�Bo��":�'d�Ϟ}O �5��`� ��b��
�z^���RD�?�5(�R��A���l����n0[����I
��mG/��׷n[�0��%�4�7rnt\:݇z���^��$���U��U߽ 5��o5�f�JY�٘~�brRc������y�D�A٥xĖ��HL���Bx�j��z��ǉ~x?>J^5G��U��|��bK�����Z�6�*^)�E(|��TR_.�2uy`�2ДZ��<���j���w�Ԅ&�p�4x��Z�lR&���ӻ�c�٢���R�_K��A(���B���h�J&h����AC'�+k:҅i���ޑ�UEK.(���&D"%�1�`���,5%2��"�V���Q:G��2����#]�����靷��P��_D��Ϝ���������ݴc"� U�s�N��w�(�X�M���t䞣�)�ʯ�r�_k2�h�}d'�i��ϑ��T�6�
��o����0�H��w��@0���Q%H�A&\������l+;.�1@>*���ħd!L����o36��=I���*_����x�>I��/̋F= ����iPG��0�z����?�gl� ��y ���7��xl���5�)?|��DR�{c&,�o��!�E�7�ր�9�M=�F�����\e��ё��i��}jjZ����!��A:��@0����������B�?x��3j������z�^��hz+����f�!?OCp+��ߧ��~E���k{o�j�j��A[	�Y�L�,//���� �~�3�r�l�����X<�"��L+BcQ�Y`x*x��0(s�-����N	[�j��n�Pco��z�z��馓��.��f����t����	=F~ �ź��E�X���Y���XA���^�6#N[�3HHٸT�y�1#����~{�Ow��3S��@�F�"tQ�+ON�QWO�쒊V8���%xL��dS��4�8�g/ю%�#�EpaԸB�.�g8�$�gm�NJߦѨK3�r�)�~�z�7\���!ܹ���ya� ��9g�8EG������E�^,�=K�
囯_�K��	AKݡ��6(|��0t��� ��ҡ���vS����6V)ʞg<������~��6O��Gr-Ѩ�ݝ/��+AC�#lH�̵V��h���@k ��A����*�MC�c�LIW�u27?'�A�- �g�����b�7.�J��A
Q)�.W�L����K�yOC����t��<k�n�����%9G8I��[�����`�n���a�޵�3i�6����)��ⱞ!B788�F&���C-����T�~p��������שM�����o������-R�����ۼoy���?F<�!�+K"N��h�#e��gO
C��O8hj	5�i(�T{�KM2�b%�\�d�6���Ç������(ef���"-][�ɫ.pDd)Ӑ� . ����2�;��AD�H<P�H$lF� �9�E4j�˞���~e�E����:����R���phM]�;P�š��Ni��� �Q<$KD�w�h�y�������W�3�.ֈH�'Mc`+y¬i��	�#-J�A;'���g����+��PU �{�����T<�Ŗ���=�#'��;�^�W�9�{��s4�F��Y�:"�@P:�CV�R�D4�=��)��c��/.	���9 �1\�pp0-~�F��#���!d4mP3k
����j,j���u�+Z�G3mts��Эp"'�MQ�+���DkA*�  ��=��R��C`���eҘܤ�~�����h@EJ`Z�0�����彠���+|�2�n�y��!��q���R	�SQ�e��8��H^̥MifWzE�0���J��X��L�{(���6�z��L���n��t��{��;�?z]9N˴���3r� �(U��f��岦�F^R &*��ª��h�S������|nOR#X����h2�x���@����g�2��@�\�r�*�"- ��Z�h2�(�(-���W6������/_��|���
u���A%�A6�� �=~0���T�1K4� O8�rسb�d�(M����#!=6= S� ��A�>6C��M�HYS	�	ŎTAV�~�-P�. ��%I��^�h�8�|1̘L[�����,ܣ\�E��חhz�2�́����A>���n
E=*Vd���ν|"=���:I^|��n����N��S#I��R�����}d'����Rx/�ˢ
����\7�� r�a���PJ$�!�\; <b���=��_�ť9A�Q	`�(��n)N��- �D�����a��
��!�����H�� ���,���=i����a( ����9p`��q�0������H9h��=������~���MAĀ�ÛS�T�xffN�ڑ#G��ބHmd�kד�t} �^?^C�S�td�gF"Y_��@�W���/�o�a����*z��|Oo�9To!z ���9�T)a���۔�̀��栎	�*���& 5�Q�� GZ$� �ԧ&h��$��LQ~-KF-Fs�k�8�P<�<5��1������"��	�w<U�40v���w�mN]t'�F��%G��t�Q�E��>nߓF��0]	�K�tF�ٳ��WB-�F����� � �?n~�bE�͂��$�jX���wN�#��#�kx�f Pn���x�¬i��DH�Ei��D2lT���q�1݃V�AA�R������\������M�\���%��BI�W�9��A�y���m0pf�e�;3ߠŅe�y��v����h��qJ�$�~W�;Ɛ�K (�@��O~�A�<�?���|� 1L�����F~�;�R!� �(y�A�	�����>��'խ���ء-��1z�ORoo7t�~뷞`�c���|�m:��y�ع�DTj3H��;��c��?gϾ��=J<p�z�!z��������g�T�e��T
G�����x����q�;�����DL�B�	ݴ�����eH��!���*	Ux-D�� ��8q����u�(��s���u[�@�Jۭp��N����c�%�!���k�O���h���LO�C�%r���)�+��0�P�
X ���{��!]�2P��`ܪ�טH��o��0K�eﯴQ������P	�T�J��&��t\9� �*��Ĉ^�-h	��[M�'"^��G�j����H����$��OpD�+H2 ��Ĕ���~�/fV��|��L�-o��D@�7j"������o�R�?��ՙ�J<*�ʓw���	!)�JC���a{|у!�v�g�RD,W�%�6����t�|�N�}����s����_���n�6r�Z��K��TV�	3N2�����FC�=W�ӵ��d1�FӋt����
@b ��{�����'&�����>N;��'O>$��W_zU����yiiyY���;����~�Y��1��>zJ�8�	���G���TM��a*V�}�L���N^��������nF��߫��I�='���R�d�����?����=zTƺ!"����>Es��i�k��H$`�9yU�t��/��}(�*�L��BT�ކxE;\�Hh4DD�vL-RZ=��Yù!*�w�v�7��|���4n��b�����[��m5Xz�t>�7�;���G���_�ycQ/`��hۊ��Dl�\��A���-zX�]H�@LZ�13����p��a��;)�qic�@F=@��.�-;�4��Exa�2;�l`B��IT���iRP(�{�M��|}��n�&)�� 0�Q:©7�6��Rw�g7����D[�p%��F��
eHT���5�n��(F��  �R�0U��OKr�M�D��hز`d;�B����	�XT3t�Ñ��P���#9^��HM���
$D�zy�F��%1D�$lT��[�2]T(�P�X��'�I6����ɀ|ޡ��{�Ԥt������s�3�S B�/I*�t�"��sNIuQ �{�r�R3xO,�{�;!�[Z�F�3�|c��k�
/ �E�b4 ��CC)������G���~X�Y�WV���FG�����C'2 ���5���#��A'�w������n6<�K����(���S�F�;�X����7�a �z�ZA�tI ;�Q��I������AjJ{��K���	#�zd��5Si����M�_��W=M��Hm� el����߮�n7��a���{��[��**�`��%�y�W�K7����4��Fz�`�+�a(9�իPh,�VM8Jtp�{� Z?��-��L�V���-��(� ݠ�"R�Ԡ�ތ��1�<%�o(qv�s�[�cq�8l�V��$a�]��GL�E��'�s|f��s�C��I�sc���h�zSr��� ��א))���<a�>������
���� �_�2��y�&h����\l����-Օ���UJ'��uV��h���"������S��
H�����!��;���}F@\�(l��ȹ�$=~���6����)��*�듼��2&��q̘����� XNrؠ���y����NA����Lȃ��1}(���_�5}�������Q�u�L�"A��L��4�E+\�f�;A�<pp�xźSUyCAz��K�'�'�!��X�͒L�G���?z�.t�3�m�+��8G�_���TH�絹�9y���!�c��Ssh��o�j�|Q"����ϣ%Ꚋ�����g�wG��]��&��/���� j-y�AOt+�����ޮ�����R�h�3��}����V�%k=�*l�Q#f��
�A�����8�RF��`d�����<Yd���?6F�ܽ�8J���h}�I+�U�6��&��#��}֫M)�BBFP�٫a�T&C�pDz�7R�G�����%1
`�D�Z���  @߿��M�x�H�� �{H�.B�;Ѩ�*�*O4�ɫ��`	lz���B���f�j  @I�����E�1 �x`��]B�̑����f��d��Z�R���-W �uBxy8����4:<Av$@�\���o�G���ir�2��I,=��z� �] �⪕lr�ag(��4A�{_?�|�8�N����W�Q��:|�3R���u�@i3��2Ǉ��t�K����⍣�'��W��޽�ųE�@P8��
��޿?�9s�olRQ�0��˗/�38��%��Ѓ�<n�	
��X7�~__�L���&t�6�`V����
j(<{��>�'�ox���~*F��b��a iݡ�5�G ��@E�X�T�º�2q|`�z�����mJ%�k���b����-�P����l�������i~v'W?z8�`���&�H�h�c\�������e�u��v��6m���N��F5���3��vݫ�5Sm����1�k�w6��&>lP����K)|ۅW���K�j��j�(a?��X����/a���@�.�.�£���������,%cDW�]�s�g��Ѡ�b��9�np���c�P��P@�의��a�P����-[�T\i0��8��Aٔb(�!c&kS��6T��Ą\:�u�D<�F��al*2�K�kh�Ǣ2���9V���������=����@z�C�T�O��,v�F�ħ\������3,5o�8�UBb����6\]]���P�o0���`)�W�j~��p]r۸&A~_�����XHD�R&P�'Bt��42Р��P�����%�`��0���q:v쨤��$'&vJ��.�{��#�%��@?~L�,fxя<�{�'im-�N����x�!���3R2�]��	�FntdT��;��z-! �׍�w��eY3(�b�r�(vb `�T��NW��?��q�Z)������/� �M���7H6�{5vymi�%IdÐC�u���xv'%�Wz4$N���J��'�롏	��qOq���0�[���I<�:�rňp5���Z�t�8il'��ΉZ���5�_��l��m7ʅ��?l_[����|+i�;�ܨ�k���?�{,� 3ss�����x]=f��F�e^8�X���"%�B$<O��3��)�.�S��/*�i�R:]��D���,�,�)�j1{�AC�Jx
]�� ���c*NKY|�@�*�\9oWZ�cЇ��Z|.%��{�T��@�T�(�	}��e�-4G����w4A���@�%�2xB�2<b���� s���g�H�S*��K4��j(&
�H��7���M1\��q��7�k�� \C�xH�#ol[IJ&���fzza��)��S����
�k/�E��Z�=�&���-��z���'ǛC�n�V+ْ�$˖ecl���q����<
�����f��Q�PE�)�3l�qK69H�-+�nu�}�'�3��o�u����V�����u��=g���^�����=��A�&�d�8���)�f_�+gͼ�ɼ
ߔeGA�09���W�Z�M�Z�q+��1%�s�d���d�⺔�+jmt�"<�?�B(&ڵk�G!��w�:���`=W	~���pΪ:WN���"?++��2n�=����7>�2h�|N�W�VA5	�<{��޼v���{т��w����Us�@�B���W��<��j���2M�r}�%VW��ٽ{���� ���XL8 �ؐ��[<��l@���_�����d�[����Yܩ�z���(��6_��?� v��3��3q<&?��n�5ࢊ��k�Ѵ�(�G�uWIR)����g�����bAoaD��Q��<���ۀ�v�n���ĹK�b�\j��>��ގ���-)}�	]ޙ�f��"ec�v����k��3��h��~x�	���½���l�M�"X�kw(;vMZ`鋟{B^x|*�����#����M�m���pˌ����@����>@�����ܸW,�$��[�E;
��z˾K���{�V���}�]w��*�5�@�ʪ�e��k�Ɲ�����a�Vj�
����e3N�ХK��V��R'��E'.@l�]h:�g���xT��Y[��B�� ��[�N��e}�� 7+�jUwƫ25�5*b�amU���q��w��F͸m6�rz���Kq����ԋ���³�� ��2)����;wF^<�"�*�7drn�,,�l�Fa�0�h}cŚfgTX�IBi ���GH�u�w��φ�
0�9r�՘CS=ը{�o��!�_<!������E�X ��c���"ۢ	Ɨ��]��j��k���O�?'�\����y���pG!�{�Ac�	�d��w/�j�V5��3�>o^\1�	��+�q�7�\8�:&��p��׃��2zZC-�s��Π�ʃF��5�K��
�q��Qb-�Q ���A���|�(��vl��8*P��f��Dþ�_cь��b���۝k��[�z�Et�� �rcj��7�O=��`�X<�L���D����52 ��	�vI�Q�#���j9򮽳���ɱg�șk�i�uyi���zT��sx�39�P��]�gU3j���	��wB�p�&$
�톽���tJ|�T�G��k�ov��I�6͘�h]M���-g�	}��
�s=�-�����3��,�#檈����Ʒ�n7"���)긏賊%���q�$\Ts���Xh��\3�w.X��G�ԗ7��K����G�x�e�\v\��r�Ъ;����&�����gCٷ��i�}(��O��ڢLO��V�����d�����f^�~t�:y���Y9�ܑW�v������m�Ĥ��R!)�=��i�++Kz�a)�ԵM@�UƢ�R���چ���_:q�4��~�#���<I�f����gϼ��-o1�eA= �O �g� 0Z5���]���n��2P�����ΰ��q�9{J��v�>8��qz͸�����T�����c,6d��}�2Z�a��NLLY6Й3�M8 �W]׫�~ �q�3�[XA�В��b�A���s��y}��69l"MR�w	���}�����(��5��B�7Uac��9��s�Ġ������c���g��d�ǭ?���ˁ}�\�#.���n.�°T.�����OLME�~7���n;�_u)vi�6:7EW�����S���V�Y4c�d��e�W��m���q���䏓�ұ�IR������/(趤8�����VXU��`wL*������5l���LwyΖ�#-�p=�N�y�ѱB�T&g�g����z�)�,�u,i����x!+u,���L������Ǉ��^b{��>3bu���\�ڙ�l��D5+��y_K�m��4�-@�:ܛ�o>�NSw��9���?/��x_����7�O�q��!������[o����?=tZM�M+�������=$��z����iG�����Ï�E;���O�%U|Fv�2���W�"'���|�+'䡇OHazV��y����o�t����������c�����]�dmcU����۞�)}���RA��C���dA�������/��i�d��qǝ�Ap�T�|�h��k��Y�
 G�GC���s#<�Y*Q}0-����D�� t��&�Ο?g>p�#X���#p�`� �
���b 2�ӱY:��� a�$�K橧���t> �ۅ{������-,$�c�����F�p��4�.[�f�G�%�~�h��Ӯ_o�P'��z��B���[e�r�����+���b>�KmV���"|���+�.�/��	�w���Z�UJ�6��Tj6Lt�b��&�m�L�ED�L���i�x�I�?�����d~n���0���+MӢ��@�
*�$P�6��Q�N����2IGK.>]��/�$��1VWͼ�(�W�AJ�M��FY������,Z#�R��m��$���=#��%�����ցg��{cc�,��զ������a�1=J��P���4/̜=��T7��S�.����A l �%���1�z��(�]J�6V'5xaS<h"��;w�E�����ad��y�v&oݞګ�8��{Ũ�6�r�-PJ�ɗn�@��ܕ��	�`I6V�i���W�Y�rKJe���ez6%GoR�����a�^�D�U��s�)����^iq�T&k� �r��]�ژ^�7��͖������:���g �b&��y���/���K���X;Ę���v�+����i�$賵&�M�ǻ�����E;�q`�k�Nr�'ùɶ!K��.�FCm�^FGRGVО=�U���|@��Ӻ��.p.~f�ڢ�ꫯ����V���ɉ��ħL2~2���]a�k�H�{M����\�.[�Uڢ� ��Eed�_>���%�V�{��ų`�3��C4/4P�]���Z�H�k�!��b.8��A���8_.�=>
�>A�['۹M.u����_�����v�4gXo5Ȯ��@>~~#le��v�3�BUk�yt�Z���n��O��_�ܐZ��ZR�f&�f��Yۗu���W��`��t�v����/ﱗNJ��;3��M�2��Rv*���@�q��y9K3�A�����Q����s���f�?m:U�/I���h���#��.�5�>̄e���
��ZU�Q� k˸����������%3E2=됥�����~�VW iZ�Ȍ���ZR��BO��1]��;�a�`f�gH���X�CW�7�E��J6?n\�3��	p�~�r���r��iy�)��˪Q�J�F֎a��s����48�C�Ɋ��AU(��{_��S'I�ɮ�n����	�,���7��^yӛRr~q��O� `�aX3���o7gB�٨��w������_^^�犖 pO�GZ��u�>��~�e���}��rp��Q':r��4!��W*Usq~|�� �P���-䀬gn90�<�t^#uEa)Y[Y�G3�^C����OU�#q!�s�1�cp�v�U۞�
^��j��D+f�ǢAY��qڱ��^Y)��aE�?-<8N@�f�g=x�8�q�Փ�~���=W�8��f�ql^S��O?����1R��+�ra�i����TE�
��9z�ov��.g�
����7 �u��<�����V�.�XV
	�:s(x�
Hli(@�-�;�,������M�d;Q6���)ը�UY:}R
Osوo�A!`���Z3
���U�.�֟��՗Gj﷥�OJ2H]s���S�-��1-A:#/�=o������$�@�nԤ�k.N�`�җ5�"�:�����m�5��� ʓ=���^u}�h���X6��*,]�˪�-�e7aݪ\��'�1
�d"c݃��!ㅠ"��G2޷4L��F�ן��i{!�I���UK^7�9	���nt.o�g�,����|۴�����/I��1�T�.8ݒg����'�[�V+���VCmQͩ�5&g�6w|f�^��ҒL�H��:`ַg\R@��T�`VꝄd&���t�+��c�ix=&�ku�~S�����vԹ-�#�m.S�r�76��2�GO`MO�?ˎ��6! �����uG��
Z�`_B5��M�O�o��DzzK�p�T��|���9o�cC{'�i�բ*,=kJ�ʪv�!Lp1?fk7�Zq��4�xe�X��B�K��EL��u��54����S'�ƫ��R�h��s|umc�bطl2ri��e��}�h��V�&;��:e\�dI���Aܣ����
�rO�/m����|�3�1��׼�vS꒪|W���F,O=��Y�����{��5^��܍�5z{���8~���:	� ������o��� �=ނ���y��`x1���g>Ћ����5�+�ynQM~�� ��,��Xƥ�=֎w�����Z"k���c�M�l�4�ud�J��nv@���9ť0��ڴ|�r:���AǓ� ��T�L��(��F����Y�%[8�tNbj�gҎ�	/����C��9��u�1�f�$��)�x�m7�ͪ&����~���d�t����y��uMٿ3'7�p��L�,����䡇���u9�ܒzO�"p��
�ݻ����߬mQZ��*��kY]ڔ�xY:qG��fg��}�v����a*)����KV��.�Qj2�|6m�B_���
a�(��"�p���#�t�=�:�Tk-��Y��H<ݒviE���
���w��Esm��w�j�h���jʕ����qG��k-^q\��ȩ�/*�M���%��j-�HN-��
W������jm�J��sA�o�����%�MYj��8�7˝9-�kf����5��/;EJhҸ/ΜY��}�c�}�����͍���,�����J�?�	����2�a�8Z �Moz��>�z� <2� ��'_��`\���B�9B��_|���PE��u�� 6�<(�����+�%~���f�����a�<�ܳv��$k�RW�1s4 �W��&z�*)yD������|�k_m��tm
��'��ط� �!��3��J� ��aa�sM�>��O�P�>�o|��é�gd��}v�������ַX��[XE<2뼠!�����l��1OQ>�K�0����9?c��|��/��n������X��hL%*�m)��Xf웫xRy�Ӫ��h�����%xiک�[H��_x�E�&T�+*G�[TT��{Y)��TT �f.��&H3e|{�+c���Z�(wdZ���LE})JՊ^'��{��������X��ԤjnkVl	ڍ�^'79$S�	���X���gd��ZRp�Y�C˭�M��*8��p��ΪUp�jnj6O���N�x��5T
�VQ �'U`4�$�_/F,��	��xJ��?�إ,^������s)�� b���o��|�C�mY~x*;./=�*����R.�����r����Q]P��Ky}C�sA��I9wj�u���� +�˚U�z��V?+�RU՘$R�/��~	W�BJ�ڊ%��/>"O?wB����T�%���x0�4�AA�i`��P�x�`X\_�0 a,']u�j���{�4�����&�;A������dAM�G�����������>yӽoR�l��.����L��gy��u����~���C~i�e���o���1�<{_1լ��� jb
l�rńs�5��/~Y��/���"��g��;_7�.處��Ǭ`�����~R�K��q]%K�u�����&a�U�b�����_?%��?������/�|�6\@>�hUڃ͹3�����+� 5�����S�)&;wΚ��g�gÔX�M���7���	�O,)戔���}�x�d�m���~�� yF���f�k�\G�ʰ:w;�J������M�Y�o�?�R2��_.&p�5��E��bY5Q7��=l5[ɖ��W�9wM��VJ�v��6Jߎj14Y5��TH�z�� ��Cڙ�q՜՜����>���[�v�4�r�j~XX,9WR#e�G�o|�=�*�V�:��jQ�料cϽx���Ϟ��.�Bq�R�@�'i˚u��]0������ǎu�%�ʉSg�ъ˩sUY������Hi�� VX}_x~]>s�?ˮ��L�b��˃�!$�8ˣkm�������b�0�E��C���#K3�息���RG��ڏ�?��5���HӬ&�gYC����'�߆ʠ?I[�&楶V�/=��,�9N�3���|p�:5鯭��X~���	�ꗿ.�K�r��y�Gp[�jB �3� ����Çf�;_�&zM})7%5�[���/|R^xiM��+F0�}�}�L�Ƭ���eX8��9mp�e޳g���W�χ�0		 ����T˞U�9f���>g�! A�, ������Ϙ� ����Ǟ0�tA[�'�|ڸo���ܸ��hҀ" ����A����� `~�{�cχs^}�a��ӧ��X�^�J
���_�2s����`��� �~�u�2�@V�e~c��(J5Ù�9���|��� |�:Hq���F�FQ��{�J����Sq�SI���7�J*'�u<9}wj :d�����?,���]�c�EkF�pqqV��������ae3���c�|烴�e�\���r��k�ܻwy�Q�̕\�b��	�K�v�?P��x"�3��4��L>8��O`��*�*=�[e��s���TҪch��u^
鼜[Z�U�cO��E`q�@	�d�Ƿɬ��M���SY���JP3NQ��g�UM�g.���c2����N=Wݵ+��C���˿< AW�t�*���TT�����O����D&T!җZe�|`��ѺϞY���79���^/9���)�O��A�UrֹcȬn���Ri��A� �7�m�td����[S�{���
�0��}�~�r�iT�y���u���U�n4�n�0�󝒯*�=�p�b��<%K����Z��W�SǞ���{��s�q=u^>��E�|�B�T�kc2�ZY�]��&�Z_g[A^���%y�+zƴ�Χ�Z�=�_��G�g*r���(`e藅����P���:~��������v��O[�;�3����K��K��"��uկ�=���ݳ_n<z��5qڇ?����耩>%%@�M�n4x��L����.�E[�3�]�7T�)�w�w���2r�[\,��~��vh�.�~����-���`��ϏE�� ��b��|�#�6���ڬ=���w)8���0h��T� :z�
�ǍV��G����`��)�@���T;k���KoVA�[��g��g����ƻ�s-R;e��/*�^
\a�
I��y�����s,�����?�3��u�^":�Q �Vj�4�K��s��5�+�v�a�\|��b��6{��i@���Ti��~��F5���2�h���JSqבhb,mM�Cw������LR���j��M*=�� �K'���U`N�9�\%�~�6��M�;(*h��!Omb2/�b^5�U�ϊe�r�J���U�
�2�s�~>.��K6!k����uMX�:˒�{��!���\~R>S���g�\+P!��3�-Ŭ� 	��ƙ�K�k�]ʴZ1mi�ǑHJ�RL]k�ppoR����{��8wB�sjOA���Qy�+OJe�^�k��5�yHѐM����֌��?����iu�\�{����K��UM��/*��^���̚>�O�O�ܻ�W�R���k2^�#7�ZEVyfZO����ܯ��3g��'��S�����}{�uw�i�r5��+��X��y4���)H�i�������)�>E�{z�;ޡ11���/~`@���'4�4����k+�ច�s ��SA���;33��uN�������_��O鸻l��O�d @��8 ��i{VH@aŵ��������C�Ih��D:X���zA�ɋ�~����\.?i��vڱ�d<m��_��!��W�t�	I��+�6tIy��;�; xW൶�(��ۿmn���ɟ4�ѯ�گ�s����r�"���4�mc�pM�9p��;�"$�{�6��,�����nX��i�.:gs����Z�7/�U2
����Wގ�w�\�]t1��w4�g��K�y��xo�{Ӏ�M���ۋ����w�>�я^vG��ՕD��I���W_sP�i�\[�zm� ZlMT݄}��t����j���wjà��G�����K�j%����P`LY�T�j��j���	H��[��P4i*xv,�9W%�����yY[Y�����L�\DO>���t�q��LT�]�陔jQ9}�l��2�.���H5l��ٳS���K>����7C檎�Tv>��x^�@�-�#ZN����'M�@�tJ|�V�:y⫘U��ѯ/���c'2���5'�NǨP.,�6�th�[{a)�ʤ�T��,���W�k��@��>��i2ɳO=+gT3߽[��[oP-l]J�g幧;����媫�TX�pfS5�/�h:�7�s~j\�咐m��B�{��߯�{���G��^`�( �v�n�j�>}��|�3��G~Dn��fY]^57>��5`@*&����:Blrr��u�ā�W�F�6x�U����a �T��`���7��n��)�V�Zv�ht��c�������J&/Z/�d-o��=�C=]0���\}�5�>�������Z�溜W���{��e��'UK&�7ȫoJ�89L-���Xr�01ǌ�y-���}@~�W�z-�</,��7 �=�*��b����gL�Y�\.e��0�/!��F�7�p��ɀ�j ܟz�)s�\}رhz���~�O,4x���`�πg�m�#��c]�\Ѣ���P�/m������7���ǰPR�	:����+���|��t�f������a+�RuO��~��Ơ�m�k���ⱦq��YٽwL�T�oVC9qvɚ�LM��7M]*���]�qU7� )��@ƦT��*���%67%Uդ�) g�1x"յ4�x�#Ŕ�����O��j]�&Ҳ�HIY�mݿU(�d��IɬVd���#��m�|˪	c2=��B>)�0-u���DϴqܻS�cF=`�
���� թ�����'�c�H��֢���'��]<���^��h㐿��k�:b ε@�)���V�W��ѯ���}��K^{�-R�/�_Q�(��	����U_��y���k9��Gd}�� ���K/�R�bמ����u���u���L*�\+7�z����
z�y{�-�O����Ux�KW�b|��*�l��G /`���]>8.>�&'s
�!��[�[̐� �k�����\����}о@��	����5@����d�L�7נH ���>5 Ӷ9� �w}�wɮ�{l<�=��	/�����ַ�+n{�
������Жq��,��]��-ǁ����|��1A�c�.s�dԊ�=����e�� ��{�2��o�!s����˿��C��i#8 w��4m�{@��ɳv���|��V��*��t�=����U�6���;�#�g\����໇9�^�w��T�+u���~>x�2�\�[��Y^��b����n��v?~��b��R-����_�f�v��}��g����b���iY]Z��Ʉ�z��A�����* �Ҧ�w;9zëm��9/�ͺL������.�DLM��|�&15���i�M�ʙfIj
��xAzN��/�?#�ʆ�(���9'I���-.��0��y�26�ZJ�$�rCj���z�$ӳ�.!�O-����������$&0��!��6��h��
�$I6:Ƽt�W+�Y�Ui�Aߥ4��X�dU���i��8�a��iW:�@Az���#G�QgPhz��TcMM��7hPѿ^c���y���Ӳw�U־���'��
1� ��+r�뎪�Z����C�\��Ӓ,$lL�"H�aRɞ	��M�p:8�����or�ќLε�?��/���媃�s��}�/7 �@����uFr�V@�`M��]�"dg���^��B��`���a�=A !�P@� ��@�@� �.���ٟ5n���_��f˳�暫L�G(0^��Po��/��_~�,O�]|�1r�����ع&���zgg'��>=;��U�e��pT�)=6��a�w��A]�uc�40�Ǉ/7����й�[��k�{����կ�݄/�#`��5�-�p���k��B��yX$�]�Ab�/*�w��eA��t.��	գ7�4�^�j؜v����(��"�P�W�:@�ʇu�\�^��^ъr�],ms4�y�k]*8;:��\��[*z��4��f�F`׹M�Ru�|��I�;{v2�	��q+�!	?PM3�N�/��J=)[���L'���$��6N5 �;�����á�@Q)�^Ss��)0\�(
訙�������d������A�c~Z���(5�����P��3;p`�^c�*I�fRr�uU�m��چ�*=)������A����)k���$�ʯ�s<8Y]���-{	�s����<$Bk�m���o�s�y�y[߹�⡽0��Ӎ�Z+����"�f�.t4eZ�zc�aг�����ђD:/���'���_0Z��qݏ�g�����Sr$3&'N� �_�����:��L�^-)}�pѽ����x؎I�o����y�R�g���=$�>іkn�nٻo�|��Oʳϼ O>��9r� ��� ���n������N{���pC�槐��L�=�ȣi���
�X��ұ|�
_�o|�?�{�k��
�4�4��FА��ޝ��e�
��6�V�3/&''�z%Kլղf� p��W�Fipo|�2��۱cF�)gyd\���ۄ9H�oaa�,�Ǎ���y�c�����않�\E�u����ǬP��2p�	�=r�e�2���ĸ��s8�����<7��������Q�=�,��k���<���׼��~���x�>h˼���s��J^O���,�{�ȥ���gn��o��� ���K���n�}E�C䫥r���-(���f.5��MsKآn;.y���(�١��&y��OU5ߺH�����K��I�%]ӋN7���bqLJݪL�`i'����)ˋK�&m�Nu�\IN�>�l]���K����V�"�BA�����FC_��l���5]u���֛�+_yB����qx
eJ�:��L+��I�Rj	�Y-s���n4��9OX��Oٸ���*�����O��l Y-���&7�D�-�C���M �f⅍����d��@ *�O���͐�ߓL�nXٳoZ����.AS��ٵ{R��tP
c'��}���$���s��ZO������}6a<��c����^9r˜�9�={����~]n��U�L��F*_7���̤	8�����w4B(LM�ԛ��__�ך_��/�h.��0?oeӚ� ����m���g��Ci׮�:�3���F�� � L��+�XZ'n�ޥ���w�)��H��C���?�� elXf��}��y�c���9 _���8}��j�۸hB�qX*w�y�u�]��R
�5=n��Y�sgN^�����/Y�+:c�$m�֡j�/.$,,�JF/��,�G�Jఔ����c���_���BUTHU��(ػ�P�|�ۧ#��s]�}Xo���qk!$|�'1c�`�Z���;��.?޽6����v#S��^�&��ǃ|V����Z�M6��5�+����r�(�S��B��
d�`�Ôă�u�sju1T,U�i� �\ZRa��,�2�k�tRz>}y��,��Ɏ�I��̬�֭إ��~�܊L�M�T� /�Z��咬���C��9~�Iy�����e����j�y�}|��!Q�iʬj8�����^�^�Ex�7�R���&�C�%�9�z�B���{8[)�}˛�Z�L��M�����E������9)C#)뛯?n�ɛ��w��gDE��f�2���{�")����j�'����oΨ���5�HV�`��"h�:���f��5�؀�{��Ib\�\uÍ���Ox�Ay�������w��{MЮ�z�˥��?d}����ء!�Ag�Y[��(Bb� ��0�0|�'At@�{Ǖ�6 ��?�#�Ї>h�n .�q�X����Z�>��	����B�,`�s?�s2�� ��
wR
�k��OF;n�M���Ԋ�Рo��*��\�`�k�-� ��t�����0v�F�c��ro (1����]��Cz����Gͷ���<�$[�v*�Q�aU�I?�������Z�վ�K�%�������p��w�ce�?�-�K�{�>��9D8���s@!lpC!�<
�X�Y%�����1g�\\�*h,)�=Ao@
�}=���e�$.p_\)�\1���+2x�]�O���&za��I��D��b	zZ�TZ���C�`mղ2ٌuL2_��6���LY�JZ��y\M�ͦT���JV1���N�v�iA�b>!�q*��Yڐ���d&2������1��Ci�)���(\=��u2��&Z�M�[����W�[���JCV��f1t�U���)�I	���GoA֤q��=iwu�-���5׭1Hn,%YJ�)iӤ��Ӽ�2�QHw,&22})��"c���$p���0��`5WK8��f�+�r�CK��<�܂�^�;KI�D"���P�U��3մ�z����)�\ڈ�^:~F��#r۫���s��O������8!r�y{�������e���q���qs]�5��?�����I27�s�nE@��R ؿC�Ւ�_T�~���h͜����]O�9"�l�I<IzߊZ`{-���Ru\��\{X���eiyuH��> ��6ɹ[���3��_`��&���TؒFI�'O��Y@�W �<�9~�k��6x�|�<�)���È�?1����� =8\=��RP�a�� ���}��&��{♜<��H��9/sG�
Y�o�c��Jd��AQ����z�y��8|�a����0�ާ`r�o����֣�0�;ϓ�_��=��G�{7��7p�i�Ag�Ѭ���q`��/�RY;����o嶝������S�T,I��l���+�L�*�附�VL�<^��~��2k<����r7U/�m����..����˙��ç�+�����MG-����"����s;��__�k����6b�/,���}s*&�4eSz~|J^y�z}9���Sǥ�c �	�*Uy�rÍe���v��<x蠜[(Yv z3�R������K�FfA!5��H�_5��.���q:b�eҐ�C�cVǙ�BH�R���1�\����?�ŀ'*� z�8BF4��]���p�T�&�l2�����`��EN�r��5���o�m�mI�_�<�?��<���T��r������y��H���l��qAkK$��t@R]`� )N���&��G�W�]���,/��?)�]{��Џ~����1 �����E�|���� ���X�P�
�k
��~�TP��ugО������w�" �5��o�NK)E[�~�|�_��US�ہ�h�������ڹq'���{�.�ga�=C�Pr��ƒ�=]2~v�X��9�I[��ww�}�����Q��a�|��>�!�DBxQ}kn]�X:���{����C���s�ុ��}�/�U,\.X:.��dϡn�j�a+�*�X>�7 υ�#�/��~��E`#��=�&� B����}��Әg��{>����nx�/Lm��f>��8;�>�	a�]�3�g��3�����W���ޜ]y�+��MMM�:��
į�z�.�5w@����1�n
�Ȱ����^��u��Ϝ1���2����֕ڦT��
�Qk`���"p�$�q�h�d\�/��	�)��黱�*��
�n]�;�(+I�����XFKG�Y8#ٍ�1�u��RS�/m��
$1�ߑ��=j�ª���B	��ZJ�@1ݵ:�*����W�@�k��Rq Ž����Fy!�+�TI�mu^����G�����/��vnk�F�@�.��Q\E�7e�g9w�-����2�ҡkD�v�Ѭ���Aw1�"�W�yJՒ�9-*���\�������5�v��e�A=~�k)x���H����Ȟ�����~׳� P���Ϩ�b�,)�h��=Q���\��"� �`ڻ�i�:��0O��^ZZf?�R����),���m\��0�{qѥ-��O��|��}��N�6Z:����bV���	���g|*%��F`!� 5�����
�. ��mo��cF���M5�'�}�{�5-��(�V���c�M��Z��ضs��p��@�ojH ]�hҧ�q�
C�po�G�6a��f-Q��3�(�
�p /�&,���������v��N7����Z4s����-Go0�}�e��?X���<k�����y�[�h/�v�΅Mg���6��=�-~;a�7?>�mK�x"��|EL��Nl)�����-He2�D'��~gSDR�
��k,�4�"$�� 2\��������O43��ڐ"��
���e�A�h=Z��z_�¤f"�%]��R��_�@�MIK��v�+gήآ_[=oUy)<kk'eU�IV���wdj�O���4�&e줴��X*��¢Zt��wnj�(�}�p3R)����Y�'��nR��7 @�ʲ�ֲ{����U��O)A�	��`ZXZ��RYJU�|�7��Q����P���s �����8x����3�YW]��i���0�'4^�0��Ø�GQ6W7�\��y��oS��v�LT���O�������t�M�j�4t����Q�>�h����p�&gO�7`4*}ٿ�-o�7����Q��qٳ������r���%�s��W>h�\�ʹf�N����p�q��r��� |�y|��ҕ�Ɔ����0����fi�ͯ��[L���e=�0���[��7-�=`���}�����1�O��=9�u9�ݮk*�^:q���V�jq�C����ܹ�&���}CO@���q���!1��S�Eĵ��>m9�h��2��4��9�{�<X�϶�s¹_�Vh�=�4�9}��x533i@���>`��?�3?3��{��뮾�,��</�w�a���U�kʻ����!0�mX GA�-���5�K��_�����
��d�U0������T*ue ��%c�|e{�~�٨��Pa��몥'\����N�:6A�K�t?��ƿ�Iևj��t�sE�����'��~Rն������4���ĤE��Z�\3���T�4Z����K7�����̴Z]��up�)�zp�6��ێ������s����HUb��!�z=,���ǥ&퍒t6��r�Z*c��z�^��ꅞ�et�h��eCI��2Vdr<'sSq}	D�O"�\�}�� �)�(�P��$׼;ȯk��wխ\�E��!�Ϧui�a5�IN��J�ّ�: ��ɗЦ�jz�-��4�	�(�X�w��^9��j�s�<+26?%�~�Q���
t��TX��*RUA��j�g�H�VU˧)��_)��%>vD�^O-��֎�Rd�+��[8/�|�+x�PN����/)�N�際�h�ɐ��7����=h7����]��^���W�wR5D�_WW�$PP�̀ ���=�s�<���O}�>����}�������� s��ȟ�ɟ����+�oXCw�0t�MS��_
Dj������D���������w��r�]�����������q;���\����Q���G��o�q�<��������z�I~��A�����U����j�Vg�0Ļ7 K�6�EBG����ˀK��4yH�kF�	9�F=Y\Z��WT��-&�v��!�M���W���%�y���Q���;v��.�
T�ǃ�LOL��p����������g�6�������bs��2]�tQ.|1��]�lG��+H�n����?�����W��
�������]Ns�,v�5�Sj��j��t��,�2hqXb�U�ca�Ri���j�a�5't���MSp��x�or*�/�q���MH�Q2t��*C}�qo�ᇩ)HY�s����~�T�nT*HJ��I��f��t�!�g�%�t�4�^��^5s|�jʒ%��\ȓ�^����J"5��=W��1���Z!5�c�>.;�2���Պj�j�蹫�I��h�I󁧓t��[�@M_�Z!-�ٖj�SF��Ϭ�� �����0�`�.��k����k8�PD�}`s4}��ȃʀ]�2ntLd]t:��U�;y�j��E��q���zgE�lH2�T�
�Ùx߁}f9-�<-�>��
�59r�ٱoJ�&�T����Q�9���n�U�����2
�uy�����w�7~���#7ˇ?�W�/����y��,P�Q�
����Y��
���� Ys�tR5��־�W��9�4͝��Ryc����
sĀkmmuȏ�jm� ̓�?4U��%'�0�0*_�l=��㟉�[���0<�r�OgΜ2K�q_��-c���6�~����а��G��✀�v�F;w�E�ap�6�p�p>=�qߧ�I��q�-ù\*k�x��ҍ�R�&�Z�<���EkVr��a�O2��:�� (�&�<M�ȓ�---���=c<7�F�b���1�.ڼ�Q����m �c-]�ȿI�E)	�>> ��kg���3�2_Βp�t�D������:�X:�/�
���D�����LX�������l�X&'�Fӂ`Hf�	�ъ��S�YPPKY��&͛3��q�7+68����S=�HnU�u�~V O�|1ay��@��׆���{B��n�,�R۸���'��ՒW������悜]=%+�"�T�r5�h)Y0Brjާz*(ei�����y�^GZa[�m�]�������W�S-W�u]�AK�d��I��°��"{[ ?����^y���'��Az%�껖�9_���F�h �Z*�Uk�P��Y��,�_R3�m�#1��	դΞ>)�����7:
�-y�]wwϓO= �ٽwS��E5�cj]�r�k
$�*��Ҩo��0'9�Oɴ
�Ӎ�AÎ��]�{��w8J�@��?6�� 0YG����������=@�׀/fb�Χ���.��[^�Z��؍����}�5�2�^z�+*L��g �'(����
y�+#�>���	s�J��(���M�	��8N��yW��}����$5��;�q�U�2�/~�!h��)���N�S7��� ��gAX��7K�E��p��=`��c_7�%��޵X,�g���96LYD+�����X�������U��қ�t�	؇��	����m�v�v/\��ԓ�[�����p��G�0^��Zq�[�:����m�;�н`_��i壟;���|�\J稛�b��������x�����o��f�E���dO���Ӎ�b��jN4�:gO%�X�j=])�Ϋio����s��R�܂���3AA�d���b 8�$n�
^n@�ۓ\�e��3/�b\�NX�~,�SM��"MO*��םۺA����XV���0R�-N�����*�5+���KZ�&�d^�+P`OgcVb�T3�߬�A"��	x9�+��l�V̯���D<f�V}���%Q.\l��|�V!��]��3Ӝ��ɠ��u{�1�:�l��MƂ^Y�h�JɲN6U�.�ͨ ��~�iw7ev>'o��f���-�7N��fGN�X�'�O�s[�陜�?ԓ�v[����WZ
����-�J]���2�oZ굎�6�����|ϻg������7�4��w��N��u�]+���_��!��o3�: J^�'>�!'
���O��#�<j�<|�%�`_4����}	�r-r���3s����Dh�[��:�'`��?����ST�Y'��s�/��G.;��|(����D绷���6�'N�x�8���nv�p��~�.Aeb�E�|0����GO|��3���RBؑ:�x(�:r�u�)P{���Ǡ�3�_���,� �`�Ēb$�i��>���!*aQ�a<w��l��
�rfm��պ�s���h��v>���nF�����G���=~ۢ��P�|���5��4S�L��hl�t��ImGJ��®.�	I���%���%�Z?fY1j��X�̛���Ƃ��H�Ъ6ui)�u�@��wEB2���ѢK��D����Ը���2=�Wp�)��eq�,�j���j��sr���e�y]��x��-Y;ӑ�).���ͳcdɨy��+�դ� �&�C��D�x�I�l���@*�m>0-{p�#�I���o�;�u"���E�����:���1�o�͋�z��O�S�+�:9�4�'����/ȗ�u]�'c��������'��[��7��m���/r������~Nn�q����WJ�\����BI>����Kɉ�M��y��*y���*Tw�? �}�	��#/�f�-_�iI%�r�+nUX3w
[�x�aO�9^�'����7�`�{*O��_�s���{b,�m��l���[�;����{����h�h��h 22�p/�/`@y��{�]�*c ��y��8�T����/�3�n`ݶ,�,������̳O��=;���-��q�5V�y��^����*J��<��h��d�-۾Go<b1�Q,�����{��5��� \�n�(� ����O۵���~��z��J�?·�Żx�;����j�q�/g�խ�.�1�oւ�'l�q8�px]���h��������;���/wͨ�g�'���M��a��#���@~~b��I�Zz�^�� �X�i_��r&K���̿k�<,o,ZA�^����N�X���ek���D�.��-C˱X�s�؍-&��_�Xj-���+nMu�����	k�/��\R��+�V�>hIZ�k��֯�n7(ʹ���3�P-��/���ky}��R]ݔͥ����]r��G���qcY�*yb}|�1��jE�K��E�«�&2.�FM�E�c��	����o.;å�Ŭ�!y̮bu��u�a�5\����K��w�>�j�8���tO�'�vK_t׈�l��~���O�U��ݱ���y\PS����sS��~jYv͟��[��/�ޫR�����ɪ
����Dv̹�`N�O+)��J��2��cO��c&�����5�/4f��y�26���������as� (���c/`�����Uc��ھ����9���<l�dr�>��|�,�����|\}`n���q��#�ՠ�
��O��O�}@����dca!0hNML�s!(�G��c��C,���umд-߃�����(�7R,�o�#?��A��N��s�p��)���+��w�ct�2WY"fM?�ޥ�n�}����50�l��c=���g�����b�����58�z{ �������۹E.U<5�n���.x���ؑsE����n'��+˓�+·�|'����L/��x�vZ�C��X^��%��Y�(�$�'��W���U� �9�����������g��i;��G�j��5����VI15�dQMW�128
�H(lJI��:SUml��;��$�ɞ��"q_5m2u�2uѡ�DZ��y��	dA���
������Zk�@�,:8�<��9e�٤	�J��mF��7թ�i��wo�LH��P����C�k�Ikp�F�Lf|�����1Q&Sm�O��u"�z�ٽoZ��^'T��w�kJ���kh|�c񚬫6W�Ö�K���Pf&�X tlzR-��q�'�⤼�w�+_S�l~\v�>(�􄍇����ΞgÃ@�k��y� (���N �@�8�K ��ϵ��倣�{�*�@h����=�9�v�A�l���m�^j�^�56&�!�55�kQjӧ[��u�r��<���34�EƐ�y�֊���X�/q��;�-�kc��b%0D:~l8���'���;0D�.���n{�p���|4^�AQoA��g����-�v�j�t��.�a�V5�0pB��X8w�,�e�n�x�Ć���L��F}�nm$�vz%xu���ฝ��;����(�G����Q|����V0����[��k�ۊ��fB�4h��ң).t����
��;�?f���q57����	Ӂ��w�-�j�)#8K��U+�tB6r=�-�`���;)�ʣ 4@�� ��"#�c�rvt��	�EPusL�r�x^�=�i}ahA�:�p��'��RP��ۨ[�E9���FY��5�L&[�̇�6T}���q�w�>�� �0�_]���%3p9��U㟳��\P �>���B����(���� \��΀�2f�����^�@��9m�)�X��.�Y����b��X�VyFz����Q�LO�N��9��f��������p�A�V.�&XP�rySn�j=��}��Τ�jl����	�y@aCcE�n��s�X5�`_~|! ���}���u���u{���|�0��<��7��e� ���e,�9�/��t��Y�.BF�V�������u�m��d����� U�W�:.��p?_Ca"2�3�e�[��]�|��sO~�������o,>g�^�6 P�d	�q��Y�:{�,o���s]_$染���>T�"�;� }g�~�~��;G�+ ���o�͏�h����v��<�q� �������\�K������l6P$ҩ��+��P"e%�X^cE��X�J�d"g�V�OH
���c�g���j�)-���-wH���G\=�lZ��	o�ejbR��j\�T��N��1�X>!aS_�j�8v m�V=�ir��*`�6�&0�JJe���\�q�q�z�\F\s�1�t�M��5!��Vk~�/�#�y�G\��V�O�3����z���7h�-|�C��R���xk\����L�H�Z .�T�}C��Z�
4�?����T�6��s��#=��I�>�c_�8i�ɴ��p�:\������֗��c�0!��cF��VZ몆�k�p�X�rEj6^׺�5(�L�t/�+�k�ڃ&�>G�gV��J�f�C��.��]�F|��wg "<}֍���� ���8?@��h���L����ك5��
^��v�r�����:�l=��^`Ϡ�8�8J�΅���V>��������	�-�����36�㳛��9��u�bq�q�����;�,86*�<xy��c/�{���v����������^�X�R@9��v��+��o�T]l���7\�~.��y����<a��K����SO=uك�'�HY�������x:.�z۴��yR ��`��Ba�4"2_�/�&^s�FY�ݏк:���Em��j�p�dYX/������L휔�n�o������J��Q�*�p2�ҰL2nl�ݞZ-|ͪ�`h���ʏKN������ZXֱ�U?�Z{^�
Zu= LǬx�$�t>o���^R- ���i>ҵ�x�������H� Ұ r0\(nb}�V(n���z���6·xo�i7@����yz��꺊פ��I�b���M ����zx�ɢ���լ�������_
,??N ]-��j:�a�jT��9rż�sc����g��Sw�&m�44�t/Lղ<ذy���]48zl�������7��`���ި�&� ��K�lQWBTG_H�zm��֋'C�w��� �5^���v�E������$�[d��s�m�L������5rO7��ӥ���m4����2i��w�Us�[T�u#���F�:��_�q��g���9���G?zY׃�DA�o4:q� ��C;@˨W�eBO8q��S�Ν]Q�h��%��BB
��${4����т�13�ۨ��;-���QQ���N+ص�w칅3�������(݂;Z-�b�c^_r��$�چ��8k2S��%jRm�rʫ�Y��^X�/~]
2)�I�R0/Ŵ�C�'�jŘ+�섔+m 7T �]}X-躆"
�tf�Ա��]������0�`k����.f�����#��DL�B>��5 �mY=8�qR�x��1���.��
�\6e��-�X�}߂��8}�:��ꩥT��X\kMŲ
�u�ӝcj�N�e��5�:�r��sˣ�z�Й�Gۯ�jL���`�]p.�~������}�����%�����B�0��,����,ŷ2�HH� ����1��`������[0{�����~��܅`�ݳۻ&�V=������B���hk��@�܌�C�v?��@����l�c�>��\D���G��vMģc�n�ب�����+��[�^��r���)F��c�G�6�$�b��c6o]lо)�������,���B/fs��'�S�*ȓY�5 ���5���o�L��a U��-S��R�o��"]o�2R
\��w���hIV2K��mW8��F	t
*N���TQΜ*��S l.+5Z��{'�K�&q!0����y犍V�����Nu�kJ*70[�%�֞�k���n��z�r�c�w��8X�ݪ�؇a�]�eׇ��ُ���Y�!�3�% ��ƚiձxO-����,M�zBr��z�<k�:��2�k��]O��jW�\=�5+F�����Fm�}P؃k�Cjm2n�� �IS��J��R�6����]<>tM�����`�Ɯ��ʨf��}��|���K�ߍ��^�x`�@�;CE]=�NFQMK#��V5^L�j���0jEX�Ӻ_��0*�|L(:^�F-��@w��_p�K]�smr������ۨл�����Q��u���cW��;^�h�2� �/|q���s�e��-`�L�V"_�nJ�V���{�\n*�,H����
�pǷ�1E@������AX]���/H�^�иqj������
�Ɏun*U �e��Z���Z-@#c��_[�*������Y9{
���LL�Ky�.�
MH/>�xz]5X�\�lR��l�����q}���{o�
J�ek���Es�����D�f�e�q���*d�*8��`ש�]��.�!2t��!x����\ϑ��-כ:��Z��$�j�I/(I�[�b�0����=E�"N+F=7� �Z\�����U3S{ц�?�JJ2�tox߾-
d���p���@�}��m4�8���uD5^[؃ �O���u�D�~��qx�f���z߾OO�f�?.*t|����?>8:�y�^�n��ײ�X����/��G��w"�����+	l^�y�u��߯	��E�\"sq�c�����_��o׶�kp�y�
�*,�*����T�\�|�o�k�鹉x����T�m+Hg�q��Q�
9tմ�Od���T{2=�C�$/gϜ6�u��<�E96 �"�
U ���ۏ�Z���N,Ǚ�u�׫�����������T��K2�^,��@�E�l`'�$<t���%�r��n�_�0Y���s25��&�;&����Vu���zF����!u)̎�X��ZҨvd~n�
Պæ�Az;	���Ik�8�ߎ�:T����w�d���V�Л��3����&3:�~$�%hX􌵴#K��NM�
E:r��5���>���=�J���Θe����r2v:X�^;bB=���#�e����f�	}r70�0�3!a�T�F���̓4�v��G]	��9����{M�b/��\� ר;!z./T��#�y4&���n��wE���v�Q���������m��ɥ���A4f���
��論4z���)/,��V�G��������@��u1 ��q�?��>o����t:OT��Q��\�4�|&N�j�?81�z�9.�
M%?W�� ��ZI���#c�l@\(��h�Ŷ��H��Ӏ|.��̧%���Vz��4���f�%��X�O�ғ\JM�Ę��Ѧ�b�m`���^�������ܔ�tZ��Sj9����K�ړ����T �y[_�Fm��!�´ڡ�[Z�\>i����̌OH�	їZ A���L�']J(�>�ӴM���E��8��P����o ���DJ�v�1�eb�O\ P7(�#L���/�A���[�ʙ{����<��Y�i2�]#�(Њp�5�	)�:�D�u ��M��#U2�ւ��5s���@��؃"P�h*p�m���?x4�7�a�X*���
�ї'����K�Y � �Ϥ�^?�I�`��p`��������9�.�Q0��
�(({�����L��nN�zm}�[}�������¨5u������/���}�>l�:�>�~~�����(��m��}����V���h|�/��w<Q��z�ת�z� 턮[PN5�4~[�$�	B
d��R��V��z��Z����iv�5�
L�j�R/��Ћe�)�O䍋�]�4S���lO���l�����)J��&qX5��*��좚}ט,3���g�����T�*��3��:@�dЖcR����ҪUp+��v3TkU0�Qx��F�ڶ�Pc�����$fMGTШ� ��N�2ӎ㲴Z��ͺ+xb��\˖�֨w�������#�X�~�J��� �Ē/@�h�]ˬ	q�)p�\p;i��1+�'���t��nѸ�1ʹcs@m�;q�Q��TaM�F�t��E�5�mu�#��4~�=h��L��i6����0G5�(��}�Y0�ڞ�p�������Ϳ=�?>�*�Q������9꫏~ƶ��h��c�f$�\�����G�¿/�ѹ���\�d[�t1��R��b�v
���b�dt}F7�]���5�;b�����@5�T�Ռ�=��	�7���;tnB��8� +FLB|7Lȱ�V�O|n2i~x�N�]})�-�W�[�W��PMoC5��R��x{�&Y��L�c�=�ֻ��}A� �i���`�@�d�3Mz����� �#�dƑHJ36áhC�1�h����Z[V���?�㙞�F֭0��ne�r"���ϯQI�j�<������윾��c�����V�P(%k��C>�읒�k���ߦ�w�t|���^MW,�l(E:�Q�2H�����+5�|��C���NK<�9[-W��bMv����{]
X[�-)R�y� |9]��\���i&\MB� +��r�JHȤ�ր%�x*�|�DO�P����GU��;ͳS_S�H�qT��t_���Tisd� G��S�k7�D\68�]/��IΟh�Y�bM�"�Rx���	2�Dz���� ���8��z^���m���@�ߵ�M���m�����P�Q��6�M׉?o7���zo�&���l�{�<Rzy8�`�@�s���Fpص̥�9�u�iv��4�`��is��"��[mm.��Œ�s1vWY,h��Kɦ��v<|���@���5�6q��P/Vzα6YoL8)����gE�hL3��"��J�b�ty�u���dfi?R�n��L8�]Q��'G��3�v��&�������z��������k�ß\���}
z���z0m���%���N�4cM��V�������S���&��`��m�.��;��/Zyr=g��A�����+�G_��]�ْP��q-4=t@iHDJ'*T���d�d��)���<M+Cs��4�h�Z9�[�Oi��F\9i�;�$.���|��Q�'�`ie��A'�T�l�L�#�BК���d���ί�a�ﶖ�C/Z>��ȵ���N�<�v���oZ���n���Z�mϽ0����i�?϶o�m����[�><nr��Y��8�)�.g��M��tӶ{�Y�����8۞��������������
�Ղ�E�M����2iw߻������G����j�\,�o7GZC������������,��O�s�s9蓰NB�W��9�`@k���'���D#lT 4�Љ	�VTG���>f3��eAh�|��PbV5�r���)�`�lX�KVȵ������EEO���},)��Z��ykL�~"՝�r���^��]1�Y����-8h!�$
�Q(�pa,�@��4K�l�K���.�4�EfO�f�^�Hb"��à�|�f�U���gy����6��3�ba&���R-@�tѥB{,%�.� 9����i�s���"@�����~0���sn1���r��W�@�}=����,��q@:޼er[���\?�v�{�}��}�b�5t��ؼ����b>>q!�/����΃�Yfv����q���μ0O�9-jP����K��Uv��H����L�*��*WK�`V��Ϡ�U�.S%���~���QP����/1�����g����=-�?����~���������b	��K���X�����:�+-$0����F����H:OݽO��O��r�ĚN��;<�ސ5�)n$�\�u�*��ctuʂO ��$L���G8\ȴm�C�)���e�Z>( ��贅�"	�Ν"IC��M N8[������m�L�mW�iĺ�^��M�v����,�l�KBT!����i�Mc?V�M%>���v�����n2��9�}�z�.�׏o� �ϳo��;��<MC|]?�8V��c��_�;�wͶ�M��/L|o��L����O�nx�f׋���es~~~�ŒϒE�F~�ĺ],g���X���Q�@�Ћ�+�?��/������3ɮY3�J��ti)@���x¿�j)km�/�ĨG5������y���ӻ����|g�;�v���>_�p��Y^��pL���fW/,�y�]Px��P�wLo��6={�
�H2��.���O=�R�ir�ї�hU#������ ݪɫ?>�n�[jOEW����`^#2#�U �Ec����j�hμ�.�44	/�&��!:Q��J��j�{&BcK�Ф��
�D���3�]i�iE�*9�x�(�ʕ���V�u���k�&��E�'�f�aѷ�~V�����������&��g�����E
7��ь��������u㢳6!��WY'1`�j�����y�8��;�1��`������Q���]�A&�Q��V���O��ǓY=�g�����c�^��w���ñ�~�5�ɩ 7� K�H�A��মX��Rr��@��C�ATe�Q`�D�ӪA$T큹�Tz=_PL�y��#�'���飒~����O�^��[��?1�d>��jqMlt����S���7��/���O�4�w��@�23p#w���ݻsB_��P3v�l�̟	xw�ZF�7��QR-�]�Mj�qC�����??04:[%(�!�7�6.��^�T�&�l��7�p� ��ϪDm� P+DY��2���^��,�0�y���XK�7��z�K�&�.��7�v�"r� �4�}�3vɘ��ma���}�ۧſ�Z���m�t��j�} �O��*�-�����i�m�h�����l�����Ms֏�6?�=��~��8������z @�z]�K��ۧP�{y�Ը�r��3)�Aj#/yt������+*Y�=?�ɠ�կ��U1AE+��X#J����'�B;t~��)
4�^�6�jШ��q�ܣqN��D�;�u�iI�Kd���7���ǔ�?���2�-�	�:#�eS�{A�w�F�JЯX�_�*i�=�/���R�	.���#[�Z:�Y_@�A֋�k�s#�T#�c�cB�<��u:�̛�(����x_UYk�k��&�ϯe�8��
�t���R�~L�01����B�vv�,21�d��\oæ ���������S���C���!,�,8�0n1H�W���A�����5����1��ڎ�	����k�jL�(wG<���Y�{7�c<'т�Uq�������o�߾��l���*kn�e�k�ؼ�ݔ%,>�� Vu}=�3�_����[�(�'� ]���j9��u�)����!��ғ�?���弖|u�v-���l��!fm\�Khd�$��t4`m>�nM������F��-\	��A����L&l0 wгuJ���;	��q��i|:�O>{N���`�2P���(��&qOQz>9���C���^�p�dl��q�B���3/εx�,�a���I�%@��!�5�>e-�3���.���TB�J��eN%�2g��x���<��4S �R�AA�E��م1Hr���r��5xY���EST\I�%H*haU�PiԟZSh��Vu������mZ�n`�fs��UA�6Z����C��i���I���6��~���|[!����i����m[@׮w��j{�;��}��a���|q~�gCm�Û ��c�E�ks@�����rX&úJ�Y���D(&B���I|�u����G�4�%t�⚅ �lJt8��x2��X�`�*ɒX�s��	k�5P$R}��b��R���hDc~y�����Z��Ɠ�:�����!AԜ�I�~�Oh� ���S�.*�u;Ҧ���Y�d�����\E����R2|N^P=k$��%¤ߥ�ݣ����?��>�tJ�U*ոĂZtՄ�B�]�#����� |`u��~q���+�����[�$�ւ+D�����x�S��A���}�5�O����	�O& ,���٦��֟S�W�Ӭ�(�|�6�L����]��I��I��&��]n�')�!�@���mQ���M���םcǵ�a���&(c0�i<q��W��j{켐7��{�?P�������?�����R�����)_�����~U!��5p���ߞ����}W��ٺ��{V����$^d�b��a>�;�s~p�K'�x���JT5y���ǀ�sƽT8ؿx�����g
`X%��~ޕ��k��i�Ȓ鳆�(�c��`��惮Ի����ˢ��r�-���� i���t�ޝÊ�>��e5�c>�
����`HI�b'��&��+�،�!�j�Cˈf�9]?��1����bc�-b჆�+^�7^������I���(uARD�p��
z�˕|�F�]�����@#�ؗ�#�t���s�n* JR/��C V�7!#!B;�m*��n�H����[�'L��"���J|��X��ͺQZeX?k1����:��\���e�/s��-��G;���h�۾o;Ώg߹�Y~1��Z7]�Un�W�	��.���mBރQ<F;�MB**�qv�}�Xp|�9bB�c��P���ߵ}��w�����X��gVE����di��;������k�G�4k��`~=�i!)�h\sp�*�}��'R-
��,e@���:$=�b!��}烌NG]���zI�˵���5]��(d{�[ԲXi�eW;*-mg�Y��4��8���⼤i��%QP�tŇ~�~�P���U�GeXѥG�*��Iɠ^�����E"��ƇC#O�~����_�י��~,��2�`�%!$�vV�������5���%T�ۉ]K_صvl$�J�WH��-A��:t��������΍�e$��,��d��T�J;B�~*������
��2h3I���d�yO-`�}�fo�����v����4���mƴ���lm�#v�����y�u����m��>k�m�_�>_5�����߫��,���惭�E)�ڵ�|3����
^��r�[|j���Q���5�|<�F]ӛo�Ѓ����.Lzz��3M��'�J֬�����l�(�O�9�Z�5��9k�s�D�\)*��Z���$��`"��&<�
�%��K֞k�dm���_�0A�NJ�	�}�օ\7:���a�gO���tJϞ����)��`Aw�h����>u�����@���hN�fcmfQ��<|(̜�"r��Yu����R�S�"�T�f�&Q�$y���W�;��(�4�U�����8X�wMB��<m]�^��[:6�)X k1X'p�w��u��J7��q�:�l���U�����k�����l����g��_�c�8��}�ۧu����k�7���nڞ��(����1�ś�d���MǶ��}��ߧ�;��>�����
�����r�>Gw�[n�bu}0��}�\�EW��A�{�
���j:��٬�Ū�Zd &�WҚ\7��A��%��Aqq̀LR�)��y�]p��J��J98�䀵�#��=��O>]�7�5隞��6x~QS�}�F�1� $+� 
�ܟ�_З�Y�_������൒�����V3�W[�'l��M�<y��<v�,�FN�f� �$��Q�����\�/Ch��GV)?�cJ�խ�H~<��EД���d�a�e������Q�B �@Aw�L
��T�V?h�(���A�?IɊjB�@�Mę4`�;=}0Q����=!0P7*س�EË�M�c�_�z��Elm�l�}ckۧM�l@_U`x��-'-��J������j�����'Ss�w_�����&�:]?�7Y�m�����VAe���~��A|����3��b˻�l��6wz����m��������i%�4Gtt�ӳg3H)Z���� F*����M�o���vx'�
�Y#�Q�Y6��Z�K��!�4�xP޲*9[�ì���/u�$�D�b�h��4�����3��ƭ?�%��ԕ�@�?{�AJ�O�ν�`3�(9�h�%������%8�U/�uo$(��˅[���J`����npg$�:D�V�TST��#����R׼"1�>���6�]P��=�ØC6�.�x�4�՝��-�,�	?���  ��IDATN
��F]4"�$�$O^��)�]_h���|���m��W-�}.����c��*�m��8{�UZo ޤ�����>Wɾgr��_�M��]ӟێ�d`���W=�}�[��~�mB�?��F�~�'���ǁ�Mo�$�T�KJq����`�o���{yu۹ace1;�[�������q*t��5�tz瘮���	v/x x2�.g����@�5+ ֩�-�J/�T9-�K)��L�  @߿n�j��0mX�$|�2]Ҭ8������=J�5������s .Qu|����8�&���K{ l+ �z���K��%k�}>߂��1�Y �p$ƀ����%���_(^��_�$d�#�U�	�5�u%�#�7H� ؽ.V���aW �<
�d���D5�fV���A%+K��y���j���7���^��d�D�{N��LB� m���ŃΡI� ���&@�����l����@s;���V ���W�MZ_�6{��(�g�j{՘ڞ�>^�}�n���'x�m�3h�������)��6s3>޿�}o'e��Mի�������|��
���ruT�瓦X&��{�Q�8�X��B�#嚐G�����>��AG�E���R���Xج�6�1W��j%��h!�U�	�3ּG���������	�܄��+:S%X0�K6-��V��`��Abc�N�>�3vEcFb�~�|��n��}4q�_&鐞]�%��% ;�� 5�%�tJ� �ސ�;��2�^�ϊ��\�p&��� �v��k��� #��BL �t�0�T]�R)�
��p4�p��$�f���4�v���i�ՙ�ࣁ>�be�hz,(��uME���2*��UrT1��E�OS�Y�WV��i�����\mn���۰+�ǷY4m.�o:�ۏu��S8�m߳�5��^ڞվ�@��%b����y���<��}��gq�t|��ޥm�c�+�c�0�|�8
D��j����P?�$�`U��N�ޡ�AJE�
/f,y�Gz��\�㭦��u#-�`@u:z5_�ߠ�]���(�Ѐ;P_�I��Y�"4���?�/V�O�$1 x��$�a�O墦��gB�uyyA+d�� '��bzE'''�)��T�=~��O����)W�5/i��G�����t���nP����%�AH& >��M�8�r�f��0���P$�SR��m'�ANK>7
���JRPq�}޿�_Q�9(M�Q�Ԣ%?�nj]������tɶA�,��F����߭��E�('<�V렩7#��7��u���#�\�}u;�Y5���d}�GȅE��I����ѫ@5,�e�n��)v�i��~���}n��iB�w��2^辵����>wM���������B�}`?��ƴo�ϴ��)��i��5�g>��&��Ƹ��x�ձ��m��~��B2~�7	�Xp�y%�3G��R,pJ���hsV#Bd�?�u�����A~���5�^;w�����Y��є���yF�5�	k�C��zBO~zN���V��M$@�Ŝ���<�ǣ9�r�9�%\���JYTR%���֬%"S�P{?K�t���R���AZ�"6ӮQ��;���&�r#��(��*��I��[��Q�	��1 EW3t�������Q�ThOm�"�W�j���S��J^,�؅�� ��-<�=�yG)�}�gK��`��__
�O�O��`M_����i�<zG��zBV�����F��2u�l7?�k,�4.����/��N�P���m>�����ɕ^�6pާZ􅭭�R<������gN�uv��_�fЎ�WгOk��p����B�����Wm^���Ag��>�n���?CۿM�5����N_��{^�6_���:f)�	���qۜ�ǹ�PE��}�{����;K�<��vC�U�W�HƊ�틡x��f��a7���M�^c%�A�3�a�"�>=X�鯿���1X-�W���x��^��Tb���+�5z(��(sd��B08)�I$KC����M�Svg��Y*�P�,�bE�`��#���E��oQ8��C�Y��"���,H�������O|8|��fEW=�G>��w�.H��*��]�2~��'�TШc]P�)���%�Hy#c��],�l4W	Fy�4�y���%�xoT#��o$�Z�����e�I���m_H�de�@\0>Q�x<:��?�c	��6�ֹ��u X����xr�o�߾Ee��$O~�k�f�M��o���/�8����^br�ۺb-p�&��q��	��,�6ٶ�=�X�������]�������~�g�?o{�^h����?�8;����8�{d�e��w���-7� �-����7>��w$9�'�����YM�I�~�EB�ٌ��9�i}V�bw�`yD�b�Z�@\!gӥ�6����}{J ��lE�4AJd6��:R�þ'�`�M^Otxx��R74_��Яt�Bf8��n�Ѡ�`�R-��A��,�X���9�N�i5$�X"�XcZ�Ra	�&"�P�W��e���S�)�>�3����,fďD�{ ]ҫ���	��+�`g�ؤ(���i�6�4N���Ȥ�G�qӐ�A2F���J��{��5��w�~t�Y�T��dE��a	���\}�a�/��~���L<�c��:~��Ͻ��v|R��Ͽ��dзY7����O��b�?�}��'D�g�t��ۄ�My�~��
��Y�ض�o�@��c�~���,��Z���A����Dm�2�p�n�*]�zx8ۼIX����q>�|����VV���b�x��M>:����S�ﲉ�����}r��z�����oӧ?���;��ɜ����g��9���%��P���?��J9��f��<�u�
n�DOQZͯ)g�����ɄA���������L�ɧ�2�/��b���P�!q�d�����]/IUd�:�[����G��G�ci���J)�9�5K�Yt�U�l��5�tL>ϐ��J��'4U��j���b��z��;�����/����:��B`��	��H+�{��LH���?@y�IL-��&D-G��C�@P-X�����M�+E�.�B+�Fᖰb��+	.'!CGL4�T���YF��dc���Izj6���>�3^��c�r�B�5��x����t����i��Xڴ�6�=���o���X�i�����]~|��K�����������ge�,m�g�n;Ͼsؘڬ�6:�WY7�3��>����?�x�{[XC vh�xp����{�F�N��޽[q����(������1�'�l��7�10���PY ���������M����F�_<���1=8�KW��p��Zr�y ���3���K�
����z%ʯ���JԬ%�
�������F4��J�B>zI�Β�nAk�4ч����+�3�o��I�\%c4 g��9�h��g`��X!$p�x�&�kѦS6 z)�bM;C�k�y��z�T脱A��<�~"���%��Őͫ�O�A�.��
��LX��{�]����#�
Nk-�BG������W�,��&%��7~�Lj��Iݦ]�l�]\A{}��?�awBM��:�u�ed1x��¥����\y-*�=h�@f��d�4�U|V��'�;f��@��e����{K�P�m;�}ޤ����w���=`��b���☄m�3��}0ٟ���m[|N?�9g)y�l��ڄ�?.�Ok���!�]!�9ub%�����v��������y{�2� �C�n�:(^:n9����~���m��5�a��ltЧ	JA;�2b�O��f찶<�0�������_�������t�������N��2�gx �b-oy=��)ҋ���X\0��W�@��V(�w8�4�B�Z���Έ5�5M@�=e��(z��+�$\>��P�	ГС�^k��n'w͂?Ȃ�ڤ/�@e�_9���D+X3��7ȅ2�k a�����9 g�/r�X�8l{]~��2-`�@�4�s���ٍ_&����C͇{E�@�A� v%M9dRP|�@�DI%[&A�@�3�p�SU2ᒈ�Q�O��vՆ�y�oJ��T�Q�T�^�E Y;�P]�vᴁY�v����6�L��gI����4���Yl��8b�{s��o|�ǎO�[�㱵r��2 ��i۷�:��3��u{��3�C�V<��{��@�����?�Ľ������w�d�E?#u��.��NRA�}Y y��OPƂݎ�<P�=z%!~v��U�+'�b���H�L8�q���%��x<n�{��^���o�g���~'�$�'G�@��<��2�:�J���]z��K�ѝ_�K����Ч���o������_��C��z��:vI,;��Q"���I��S�J3��B��0�F�.� ?�������a��׬�wX�<>���r%��ٌ�u#��C��4+�X��T��������㾸V��@�U���H'HȠ����G
�.��"�<�>?X�������Vs���J&d_8���m¦żX��*x7p�
�z�kuÐRhg�F�1#,jHt\��4�ߩ����Q�RDe.N��Ms?�q��'�4�H�$a�c�?�?�5��a�!��(�ң8��ʘN�~���ϧ�p�@b����a�&���v\le`Ӕb��k������M����'s���\7�Pn-�]���׾��U����	�}>�ت���V���_�R}72��+�_��V�\�\���X���b+�[�^�����f� t��c�-�k�y���V~�|~y9��<�GCh��]�XOh��j�)Xbv��zY�B`|Jo������^{@������g�;>f�}��z��s���I�A��,g�^N	���&~� �3�NY[�w�	��
��T�(
u�����)�4G��\;0%˕sE����$⣰K(x�a?�k���*Yh���]_:�P@�f��H��R�"��/��
��岫-{p��~�"$�,C�o����'dB�P��Y��8�h�t�.�u���+�@��2 d��_�|-LZ���xL[����@�j3Z)�B�X0�Z5g�ցEU��s��&_�b+h<�f�-*]D6'u���������C���ǵla"������x��`⵮�M` `�֧�a<">�ô2?;�i�^�ŋ=����
�r���)���U[za�i<V{������nc���&X�gm�۱>f��B�����e�	���ݯ�g�Ȯ��]ۻ��!~���6���� ���q��	� �<�8'����X���q=>��@��ke�b�|�i�O�n"Z��M��;�%h"�Z�Q1�ٺ��4�x��Nǯ?�����/�������L����Sz�FC�Ku�,f��s��z�lA���/��zG�S-��T�4ކ� 딒>	WK�7�)����<xJ4'>��I0�C��qLƚ�¥.��1J���A"4��h�� L���l� ����o"�HnR���f��8r�f��R��z 7c�FN=�ي՜z�	�h18�X���@N~���p	�#N�M�f�� ������S�[7�-Tm"�J���� � $K2u�`A��X����R�6�m>^3���ķ��޼��f	�'���>�B|m�α��c`��/j�ۂf(�5��׬�5�k��R������L��>��~_|n>_�cw�ݫ&�P��b���b�x���������]�>0G���9�Ҷ�����Ј���~nĂ�[�拷g�k8l����ߩ�9��go����?H��M�����=z�����M�B8��irr8�:Evp��Ha���MFFf[w����G�a��?|@�~�=VH��kG����IE*ASd�|qyE��kВ	�:t<�� ��w��)�|�o�{\����ݮ��#K�I�7Uf� ��I��D�#�`m-Z{7��od�@�􄓆'%�Y�&��瑴T�I)�t���I�N��"�M�X4Z���l�XP�5�ˋ3�w��hd,���-�c�p��pGI�#��i��L��E�&j^��-��-�A��D(rm4 �k�#+fR� �`UΜB3l\��X���.���9`ks�`�[����i����)vYxM׻<�y�ߏ�D|�u<�vw�V�}cm���x�1�j#hT����׶�-�D8���c����<Hڳ2����b�������e矩W�~^{A�:�	+������m�� ^I�˞�t���6�x�?~΅��3>�v�5���7���5�h}��.�҇��+��K�NSm`�{^�)#J�׌���
V9&�����=����;��?���ſ�G?zA��08��D�0��G���4!���z4�R���Z��
�_]�y#-NB� }aa
�(
B�NY��@�P}B���+-uP\U���[��\xk��lK�K"h�Zvp��W�W�|�C`��!���Y-1
�Y���6��� �I|!]�f��\�>�
�i��\י�l%�E&�T�b��A4?i��@�M��۔f����|Vi@��gP˸� �� �~#�O�}���i�R%ԡB6KsRw��Y6�����6��m����X X8V����z�}c�?���G0�b e��9b����ݧ���#8�>h���j�\bA`�ƻ�|)��,d�yv��|6����6Q,�b��k��=�l/`㠧?��բ/����ڶX��V�=Ko��l���ޅ煯���W�dK�a��,D�w9g&M��໿����ko�����):o��)���ǴFO��OZ��`P��;n%��z}�m�y�i1_K���ߥo�ބz�v��k��?~��j!9���I����c���ܒ�,3�u]Kja��B�#_��e�8D+^-S�� /�P'�M�4�~?�&���Ч/ �m���#i���y�k�C⼗���"��36-WM�
U�E��E�����{�'c���-����as^XC�{"T�B	��xr�}��D��0�j��o��2�2���#^��u��6@�e�%��ڷ=hZ��HN��ɛ {�H�+���ikB��lM�96R������dkY�B��l��A� �&��}�F�5u�	�ph��&-ʳ�i�{��� ��G��;7�7����~_2����2������1^;�=�X��c����c�?��������������-q>l��>�'���2����5�s�+~�ٻ���7�6�q�A�������� �dL7l���}@�}����g�gp����⊎�Ҫ(E��i:+M��CNv�B.�5j(��<���������u������ӟ~LǇ'49��g��D����C�F��֡nfK&t��DQ ����@��`-��]#�OL�Ryٻ�8m�w�$K�b��Zs&�� ?�=��=�䕖%�m�'�^��ʫQ���$`�����5�/sqk�e�rI�!u�dcl��������v�M R�V���S����	. �D� 69�M�l�>%���zCU�%N�WKFA9��*�T�h	�	\?�N��h�"��H�F�(����@�/Z?��D�n��c��/4�Q���c�ͷ�����ۛ�r��a��k�]�Po�)�i�8���Իpl!���3ނ�6��*K[�q�㴸E�L��a�c�1��ݳ�����N�ޯv�u#ٵ�������۾���;�\6�����~\v����\�~�������K^���^�y��1��h
,�[��/�d�ϔ1��_#M}X���O������1��Ǽ�y��=��@'4����l�D�� H�����<��5Q�XBSE���iv������<Xs?8����-��GO��`0��x�!���:@�,Q-:���nx��M��^�A�신M�6�H��#�g�Ɏ�)�%��f�P��D�������x�
�p�!�2��aQ��A����T���vU�XJ� i�`;K2qK��?�������s:<�Ke,N�xB�V!�ɂ�|=_��{�V���,�Y9f�* 0M�	,�Ui�T�"��#x��:��ӓ�E
K.$�v���A2yB@W\<���4}���k�~���i�>��6[Ԟ��~{����_�t2�X�wf!x`�f׏���>�{1��w?y��>�T�XK�ӻ�{��|>o�����g� Y�h�
�����6�#�jm�&Dm_���-��k�u�؂�!�_������6?c*g���7�}x@���m�z!kk ���Z�|��5%B��>?>�s��ݣ[l��ko0�	ȃ�e8�Cw��V����{ұ�2�d��X%�"	߰ +�<B,>�� ��|�z���f8�����駴�H�.��K!�-X��m���� $��Ո�\�"��p-�g�FUf�/��R�l�}�K*tl�-��f�osB�ٲ��f�*���G�_� �;��k��s�ß'B�C� �:$q�X�t��|��L �3ՒjѢ�˲�6��Pǋ]�@�1�v���R6���q��MbiQ�-B,� �U̥H�/ L�p��qk�＠��J�]YPKT��D}I�w��/$�����>~`�4�Y�"��4Ќ��LK�k �X�b�k��-`���iZ ���v�ǻ��u��i��m�w�x���D���1MЃ�i±Ń����>�g�ׁe=Xڿ�k����ێ���}f��1{��|��m���m�?�p�^�{׌n���@7�M�ڽ�����%�=�s�SW�w�����QrK������H������6t|rB����R�����8���~DnHef�R��%q�.Ο|!@v�������ߧ�o�M�|���/?�.}�������V�5=�Hϯ��� @���j�`���qG��R�`�/���J#+�SwG���_� �h���1 iH�<i�2i�M$h�Zu-����N�jI��o�QM�e���{T���a�zU�Ͽ(4Љ����BH�4�()�4�-��2�;�a PY[� Sd9�|4�X�'uŤie= �%CH����N�iw&��obl=��]�3ZҀl��z���*�`5�P�I��L ݼ ��G��	�U��[��@�&�Ͻ;qc�D���s1�; �Z,wp�V��)v~y���g*
����pb� �hM(`���*�b6W��5�j����2��g���"��n�M���{��,?@sa,�j0��=c\����
���0FsQ,�ó�������)���ɸ��Z�s���wc�ؕ[����f_�^gﮱc��g~kw{��Uhc��!3��{����L��tآ��u_O����Dε\#lj���z�2�֢�u��uz����ݧ[l���)�)���]��´��`F����h�(��yI��恮�w.u��н	����;g�p�Zo�����޿K��}���o�������1]^O����}@ZxT��R}��Q�3a�U�[�6+�#�v�_�1�N^z�
�K��I^�HZ�;鳵�XދI�^(}��M���FeB�>44��yuyMW�s::
˜;�^�� ��9*�sB��e���E 9�f�2i����j��Z��~^f�[��!�EKn~ư2V�K��'X��5�;�f�i�j`��!ް)dJ�M��A����pU�i� )[��4I~�lљ���W76?l -�½T�OЂ��: ��J��
�� a=�s<kԆt�:;��]�k��轖����x�^��i�����z>�ڞ�����n���+0!�]'xgv{���L�pǎ3P7P d;ގ��{�ރ||��
�q;��C#M�w����ywM[L�ާ��A��A~#�C�N�8�}���dG ��'��*˻����N6�?$��<���P�N�|M�����A~� Q#��-�Mjq	�v��߼T�1�䬉������$}W��ѝ7�~3�1ȿA?�����?�����5�ȂrdZ5�z�l�4t!B�R�> n��T?
� ��t4 ��S����8�k���|���͗/���a`��)�l��Bj�<IA; �3]֌�cVS�������4��f�uC�@�����6�Sk�A5�Z$��d$4J��b��h+B 2RJu7�1n��t΂�@X�͓��4��-���4g^>iX����c�[��Y�&�2�6�E[DbP�ZCJ:�mz�v��f�u���@�ⵅds��ڙ �x��)U�V��[��9�@��T\�22���6n�Yօi�6[�^@y�Ul�x@����9�f4�k�� �p�ߍ=5��VEǆ�.ǚ@&�M�	�1u�LiB��Z�P���X���b�6�P������ݳw��8@���m3W�w�y!���v={�&c7^w�s�Ci1��ޥ	q�e�*!�n��w�^�ً�[>j�l��Ge����o��o�#|⒁�fR$�|-A~xM�F�䥥��:	)y]p��͟> %�g�暧���_�=eT(��Bd��4�C |Iã�z�k�����Nr�ܫm�j�F�e�m�\z��E؍h���Q��KϴP�6����2��H
�mo�<�E?!1	>@�O��4ѹ�<��c�g�'ݒ�y�t��ԬizU����_^�_zGH�z]���S��Uj���.%�,�_��D��3q��ģ4h�\�a�8(h���q�@s�D,`��]�b-,gl�CaO ��f�Bs�W��`q�򚢟���j�}��ѴA)�Vl���]]]m\ ����/�l��V�in�T��۲b�߀L� zd�3	K�r���U�s}5ݦWv�)x> �c�.��@��||��=H�s����KV������{�1,/ ������d�
���fɘ���m�	v{�>-�ZכX��ٻh���Z����n{F^��3�콘�d���{f>;iǍ�o��ݸ ��m.XL�[n���xb�����X���]g�3m,@)3�����C�L:ȃ/Q�4�� 3�6y��� �������Q�G������JBlh!�1��E�Ìf�Pә�4�X/���h��&��҈��X���?�Z�xm��c��W��jo� �܏
d��'�b�4|�8��:��K��������z�z��>@@���j��7�?�U��|��,ݯ��v�H�A�_�d����y�P WЕ
�k�>�u�s��^	��V/�����b��L]X [߲Zb�ۯ�t�B�.K���5IY e=�f�/0�0Vq��)#�]���HSk}�]��Ȥ�/>ǄNS�ҩ�$�@��q�ʦ���f ��.zҖ�aam3iĖRMNxy�u��.�E$���sf��Њt�	�v���f�N$����B�� �����Ѿ�ڟ	:�q�)L z��@@�Fҙ��i�wP`����q^����&P_�RA�%z>�u^�K��!�l�V����^�+qg����k$oXup�`����tJ{^��gb��sP�٥�ج�Hk��`v�X��B@������٭�n�)#��\�J,��6H.��j[$e- M��C������u�L&ؕs�ac�|���:ِ�1��T[�FwM[jB�h{X��ݻ�O�ҡ�BW-�#�%�B�b�F�����z8�uZώ�Gs����ր^�Y)t�פ6D�03�vL����%Q_1i�wxih&RC�P�t]{�;%�J���i���2��"��B��4JE@[�)��n.�K�5��^�N2
x���V�=��y���$���΄?�Ev=��g�e�$�+101�>�����W��L/nb�<�ࢂ F� ����LhΖ�tzF���4<=�E�A��TSdר�e:c�:/eD����l�=��&�I7�c��n�E0�D��e��dG�waE)��ڳ7���� ��bm�ƌ�3��i��m�^m�4���1�ǎ�2��� ?���vL(X\»r4p/����g՘0��o83/T��鎠6�b,o!Y|Þ�=G{��}N���tpp tqE�l�u��� �W�j�W���;�x{ύ��3{>����,�q�{7ܑI���M�٤�}W�n1�C/�����{��5��P�=�_��5Oʅ%&�R�y ���X5 L��ѨKF@�	�u=�Ol醢H�p���4��2��T*(�'��y�=�ռ���Gt����b=�F��Bp�� �j�O*�56�хvyҵ��Ŋ�f���@��	�#ē���s�vs�PD��y��d�/1Q�	�|y&P�3� �&�|�ke�.�̆"��:�ڧ%K�O������1�s:<0�dA�Cp�$X��	�Q!�dui0ֺ ���H���B�Z�������B���;_ђ�㲆
���ZQ��ɺ��y9�e���8�7��zk�b3�G��fߛ�o�U�%���_π��u���Yq��Y���&�� ��7U���M�:���m�����0W�?�p�g��冩� ݄��y�1d��&��jZ @�vM�m�����5i���2����Z�%�����Fx�_����Xz-�]��V6Dچ��s�`�)���M��.�e������}��rqZz��]=��{�$s��G�>n����so��~�����ڐoa���b��x<�s����vy����2�&O�%U,-�5���tDDnz~�&-��{,C�!�4��/����z-f s��%����$�>��z����w~���dJ���r�{w����M�������i��Fs�+k��sC�[6��`�l�+�����.� ���ڝ�wA\�x%�&d���p� ���r��v\/�����%[6XH��]̗`���2=���LiHՒ2��|9�wVJ-�m���$,�J&x|Lӯk��h�f%i��O�ە4e����W(�`�O7 /��9]o@���Sl=g��ϓ��{<V	
� �������{�7l@�ML8�b�y�l�_���-.<;|�gg>e�l�6-@jf�׬p$��i6��^3��&D�%#�4lo�X��i�m~]���{7�c�~��eU�>�gJ�<�a���1pmA� s�Nx��y�J�5���6�1���3���,-�m�	+�_OQ!�4���U���<�pºQ�i�5!�a� ��:�.Q��E~��8V�݅�<��m�X���"J�\;I(S�N��eU(�˵:(d n֙��6}�w���i�q'�b�?���������/�.�;�"�f-�)@���� �,U������ �"E�-�a�r)K��jA���,��j-}� �b�I�ht��ߣ���w��y��C���irW�\C"q�L]:�h��̎����"D%�|o���БJ�L�z8tBg�,�
W�z��<��41I},�
�r!�*�[ꏻ�=�\,X׸_m�s��d�_��d8�sI�6�	x��A��Zz��@ĄX�!76���> ��R�v+��%�^��.����C���MWX �Y[���*�K����j@���؃Ԥ�YK�ܤ
^�N�9uV]���O���S��ܚ�ڲ��bm��ɾ�䔿�kz޷�n��N*45d�!��a����S��X�R(�1^d����[\X�˕��S�=�����r���а�}d����@L���%N �{c/����@�=�����f�.rt
�<I��+>~8���1��}�W	�sx��˱X�#���舞�x.�X	O�?��F`�o���K2�F�%�
�߲���U�����&����]��[��9��el.�MQ��{�͆ڸ	׏���d�^���L�F� �\o������+�4@H�y����8�]�%(�
�&̃��	ϥCzŖ/���XL��������ߧ�Gu}��/i���f�:Z�0]��îfc�Q�_��*Sj�@����9��e �4�|F��X\W�3i5�\.��R7���7))�]�C\�1=A�*0I���N�*�ն�f ����3�Ǜ�I�~�@��BK|� ���"��K��Fap�`����F!�L�`k+T�G'ռ��nLE�hD`�� �Y��g���/X�U����j��.���������2!�ʉ����.�d�w�G������x&�����ًs���y���\J��~�>9͕�G��eA줖*(���yƚ�%.5�r��T2_m�?�Xkq��΁�L3�q\�gn@���1-���r�-xh`k@n���2DH�k��}�0A��7P�#�q�3㭱��=�fA`��Ͼ1�2��- �?��%�� ,M����Qx��:����k��w�b4����ZhB�K��d��X���3S&�ƧZ��7�	�*�;�?���7�&_���x���^TvoRP�\�w��[�~�/���̠%[Зg��eQyW6�G1FBP�J�\�B���g��ht��>��_�������m.i��?��w���9��'?�?��?�w�q��heĚʘ���1�t%َ5�RK���)���5o���<8%����h1�*P�e�� �f�vԬM֊hF(P*Lϟ�u�ZMY�V�F}���S"�b��B��K�ˮ�_��[�B�V������tʺ���P�hը��Cj%#��𦢂�v�	Ye8���֊Y)t���) 0��֜*q���С��h�	EMC^��<?_��g��Y��!4��Y �AS�D��V�ˏ��:���9k
 h�[!@�fHeʠ�V�%�Zmi��.8~�s�Ż������گ����\ ���]�AX�������d�M�y��%��
]��*W跻杖{y�66Ӭ} �s�[�J4@ɯO�K����`n�����ݏVԒ1dl~�#��v��`��������o�s�M�3�?��,��c�~��xA��Mh0R��J|�&�޺���7��ߣ7�&�~ru������n	pC]�i� ��x�2��⇖,�&jku�j#{��|��q��G΁^	M��b�Tg�7r�j捺\P%��梭%)�˨J�Bgi�Q���ܱMH��*����P��];&�G�㙦���7��j5�����/^��O|�ڳ��o�����]�ї�F�N�ыgs��ߣw��@|��������CY*�)[ ׬�/�g��˟��� �x�dC��4�<|�m�����)�V�l�w��#���b�jc��^,��t�e�,��jQpG�_ >�j�3j���M��j�:q�4E;�<`5϶Z���6Z<mK�,N�R7ʝS�߭`�!�Ge��+{�"��u��r�HU�C�3����W4Ͳ�k��r�fg��} �'��s�j�![F�I��Ņ4\��W��h���=��92Elm��>�xzZPF��	D�'�	�߳iU �E����«M�[�kͪ
*T��΄�r7��s�xM�ޓi>���Ub g9�����x�} �5�Xbו�&�R�B(�����X�,Λk�h�m5wӪ���k��6w,��ߟa�>��]*�X���se�w����v釁L>oQ��P��hFM��<�N������y܁�A}�_!���y�̈ĥ�� ��ڸ:�!���6��ҭ��H��$٤��`Y�"'[��mw!�T��(����C�:+��tA��Ƃ�A����t7�K!�QT���y��.-F���%e�X��ÔIa�Eh��Ϛ�X��������(%�z:���_.�� ��{t��k�s���������3؟ѣG��ɏ>����ߖ����#z��w���&��ď�������.^<ޘץ���8�:����tprJ�'����]�s�5::�#�2��ݔA~uA��3�^<������1r�%�}�(�,k���Q$��̂���_y�Fy�l4~F
�ZF���Y�W��[`���&R����sj���
b֕��J�+Ჩ��cT3T}o�.kN�J��U�B���#٭I%EezW:Y�.�bZ���4&���BF�P�׿v��~��~�!u{�t�]�`��t��ϯh�L��Ƣ��B���)�'AB��ÅF�&c���Ё+,j�0 d���F41Xx���CA�vq�!\hA�I\:"��dE�&�M��x��S*Uoj�5�$��Q8Z=RP
$�����U����$hX�  ��g�KDW���K���m�l�L�KY�x�8&di�a>�%�����۠Z��hsg@{/�>Pų��R��,�O�@Y�mǷ�J�������- |ֈU%w��� ��@y҄ �Z҄1v�h:d�g�3Z� �?�T&���
�T@������/i��l�m�*�Ư��d��ŀ�UH���Gn�y�����[C�]�����$Pp�Б�-���I���v}�8ֻ�J=(1E���� uMX�n\�!��:z�?����������m��،J�p����@?���GD��o�2MY��o���B�=�#������?�������� @��{q�')��}d�!i���:`m�/;gS�d�����x�'G�t�`�ƻo���C'w��;�J�R?_��Lh�ͩ��y�	��$Y�6�hL#O)S����	�|d�o9���ܒB��  l�M��j ��������p�,T�
�H]�j���R! �:� ���6B�XBLTT��#����]+A��0�F�(L'�JJ�*��@��Ä>{��^�8����O	�Qq>�Z���T,��k��Cq�hN��j~��pBx�խ�T�8$h�h0^$�i2�8�4�v[�AX�qSH��]�*���_~���k�Ԃ��p�[�0�s����p�S��ƴ*����I��LS�n�p]�c6����>�������mn���-���c���攅.]" �e$\8�f�!���Z��/V
��l>BH.Cj.4|�D�~j�~)x]�_~9gKh8�y��n~xYO�n[@����.�hm6n��z��:���d�t�K�^q���M���[�b�Tup#'���n����?��8�yc�O��]}��1zXU�]%���ndo��"��gs�ŋtzz*?s����~���گ����;���O���>�fI��<�99����}6���/?a�Eˌ&�����d���ՓQFNO��ٚ�WK*.���+\i�����G~-�F�G=��M#�cɠ����0�iq����o���fX���)���x�M��ʵ1G�h�F�=��Pē��Ԣ�&IMJ�X�6�K~���i��T:�6/Ѩ�7/2Q�9[ ��	:!)��Z�z�5��m��9�,������B�#��k�T~�&�����>&L�I�ߗW+���5�Z�z�t/(�}�-�ڃ���	k
1sIr��
$�`_m�	��"��d@�`B�FL�M�sYJI����'>��q5�����-t��1�� n��ŨaU���\'۪L=\Pu0�q�p|�US6�K�T�*����qp� ��q���ȇ��n0y�J��}#�j��(��W`�$��B�ǑhU�`/�Ť��n)>��jn�بxJ@�Tky�"���,�?�j��^_3}�=�e���O�_Җ��ߛ|V)�k���s��[�"��Ym�4	�U��>�}���g��_����Ҭ�M!^��qvM<7M��R7�V���e���zK���6�dp;�繸�|����ݻw�꣏>������R�k^��SoB��%O�>k�C�0]�����a�(g���!�./h}���Ռ����t2>�ًg�"�J���,V˚�YE�ۍG)={��F����^\}�W�Ui�C�ggt�a3o)V
O;r��rEk�~�� e���Kb�L��k�U���L
S������)�?AR��y-�wM��ᡠ��g�f�4.�g&��6�K�1�,�Qbn�U l%�;��`�����(�M�`V�B�B���9K���H�>M[\k�U L�\��U�����-ł!,��O��<�
I�%, Ӕ7Q��Q�q��Zd�����C,E�)B�<��~�i��;ݼ�bKw�&ǘ�\5���f	����6JS��.�/*S�Z)�{2��B;��1�e��J��H=�lư�J�7��鉺��B��ґ���[�F��;��P/�{��,��k�����^B�T�b�MM��^#YMpm!0|�
kd�������1v�
0������4ܡ�ւH�.Zc�ǌH��b�F����o��7)�u"�L�\���oTY���;�Uʑ�%jޚo�c/L|s-��U��V�)-�d�u5H[�r�l�Y"�	5Ei��J��[�ъ���dʅ�[�V��+��� v�w;#�������y�����y�X��	����wNM���9�xr�_Ni�R���w����^V���`Ěɺ�Ǐ��c�8Т�����E�Z�������u�Rү~���=�򌞾8��~�3:}�z9��௾I����s���5MNFbNw꜆��/fZ�"����:����Z�db��͵�wW�jhBM�y���w�5�XX�YQx���MѠ��4�S5^(aT��R�$�>��{Ǥ�b���J�5U �
ENkM�`l��A�T2��P����S�3��L��p*u��D����̂������� 0.ϴ�J4?��E{��������!��Z�t��|����G)��5�
�%�%����.�s��J@��<�D����c-�^���4��,V�L������<δb�Jޥ灡M�	Ne$1k�*d�����������`���Ȩ�P�~�������،�D,Y��$C�N�v���lѶ˗s���[7B�l��F�m�jy�[gJ��;H��fW�BS��>�d=����J�P�l�S/w%Z���ߎ-XL"�Cj�(�gE��@�UJh�ZK��e�PJJΙ��ĺ�0p�����o�KQM��6��v-S�)�[k@�����m
�@��ص�jw���0_��t�[Ϊ	�O?��rХ��D��[�}��-���<?{!���߷,/�Z�����Ň]������'�'��<+�4<<e�=z��..�t�����t8���/ӓ���b���Q�F�	�X۞O�����>| ~fd|�}�T�7=��G}F|#C)�?�P?-��/�r�P�����&���Rl��t�ЪO����S� �KUF14�&q�T�*'/�D��� ��h�y�������N�ג a���Ed"��^�EP|C�X4�m4�G��HR�P%܄�%�d$ckfŒV�@!�"%��N_�qtzR; ��Y%��8�{]-�d"y� ��:ݎin�N�T}��%�A��&��YB�*A��#��xV��8
�>��^�CZ��JwA-E2*�ĉ��]zgA�� 8ƴ8�A������m�ߖ{%^�z�m�r|-��_��`���ҶX��"Hij�;FS<d<�<�%�J��-q��Io�O�堟�'K��=���F�q��ע9K�*��W~�`�tm�}���__��n���cQ�%�-��@�*S�7�e�$�ρ6y�J1�O�����Z�\<?d��/��o�u����+X_�Z�um�h�݃�cn�Mb��4���F),�a��{��Y���3�jW���Ν;���� xN #.C�W>��
�[>�)���ٟ��SC^�RH���>��${�w�w~�7飏>⋬�����O~L/����qF����(=�����8��hĦ+�O�P���@���##a�����;}�>2?ƒ�vu�����/<�49�YT��4)͈�4��ǬA�|�� ,4�&d݈�^*C"���pЗ\x��%,�F{��u�.��<|�D��4�<		���TiV�j_�hf$
}�S�����>g�(���ų^�RTI�_@�Z���MSs
�$2 �i*]�\�rEh�������{jY�4�\5"�G7}��frp�HCr�u�A����3�W��� F�Q���
(P�d�Q�.�538:���V����r��s���R��L��^��[x&PR�w xÛ�t0�w���=���6���������|�5�Z�o�"i�]���u�o�i�"�~������,��qE�1{�Ea[M�]�n�˭�i1,����b�������6Y@MC�P�q� ��V���=w��ۿ�`����J�m��d��'(�F+�I�-��Fi�a�yD�3�����|�u4�`4T��@Z�<|�F6��>���vzz������}>����/��/��f>�Wtv�����+t� �DA|�7��/���G?~Do}�!I?��Z�]�/�΃�����|�����;UtL�~��J��c)����ͮ
:be��t� ԥ��3)��38�X����Q�I�i+5��C��\#�_� �,�MH�MC$�P8QRZ�.�mzH��iz��6I�]�8O
qL�/M�B��E�/5���l�Z
?��5��0k��Z��� ��p�5�q-)pkɶ��
k�~W�o˾V�������PKZ�%r���J� .ǆ�
״Y��bR ���,���v��whp8���Ң��1���>?@��e�/����3��ߦ�vh>�F8�$��{�-c�z�b���+m6��4�]�l����?���UoXE�o�i��8n $U������8P�VN�Mi���6c$4aS7X�?��m ��g�Zw>`�THI�s8-�]���P�c���::ֹ�@\ּ��Ǡ��N�����%��+�}�sf@a"f���l���~�����/~p��>8��%�f�jQ$(
5�7�p����ܩ
�pG��^���N瞳ǵ׾���k�_�I�,m���Cs�3h����
Ӿ�����)_k�%�Zr��%�;�/��?kO��9�>�g
B���Pc���������~���7|��}��Y��#v�CN�;�E���V��V�r6��������$�e;��-]���ߠ�wn������L���t�`�.�[�"i��t��U��p�P��,{{�z[n���#:?�H)?@��-s��n�UP	�� d�a��ݮj���HbYq�q�(��
>qn�l���=V� ���X�W��/B�&_2���-��G&�g�%4?�ސ":-�Hnn�v�6"����!��;�'2I�t�OÁ���,���}gi��s/��
��M��ݟqH����
��D��M ���.b�=�R\�&w�����
��UA�*$���im�U�e4<����a!��uE�5a��ۿ��A�-��+������f|��HB�Z�%T�	�zӎ�b,�_���{�Ŵ��?�Y��}^?<�v8�.���m+��d�|tsR�\��\{��e�Ϸ������Q�K5�YG����zn�Mo������m�DB���tS��Z��W�vS��(j�o�P�vE����	4��|�� �=�(�;��@�P	V^��V�e�K�(HDHgg2�!n�7�˻����ׯ���W�:�6,̏O�tr>��������w����?�_�忡�~�2�	��Y�O��勘��ѻzp��lN�&,�٪Jf�����vFk���:ػ��b�=s�IC�1�-C�F�ĩ�4�)]N��tr�	8�$a�v$���u��e�ь\ϐ�������*��\PFBF㜕�LmF"�u' ��'|(t	?�=�"u�P�-�m�2$�l)D�
��!��:s	� ݝX(/X��� ��5�Cw�\�N!J��bQ��n�p �)�v�r��+,WX.�J���c�MKH�CbG}~N�,�(��p���ꐕބLw����=9�.l�XJe�P1��í�*�:���&��ߟ$�\,�yOx�,��Ap�]V+�����t�K�z��!���5�������(�,U�ۖ�\��.8��XU��)�"�e�?��W�<r�ݢ�[�F�yu!��r������`���P��6!�U�IS����Lqu�Q%�˘xM��j]�>:*O�:�{3��reF$LQ�sb�����mBx}��<�Co^!x�ad�{��w"�B��umҭ�ˊu��=d4r�����!��s�=[�4������	�iڟN��=~�oy���/_��h	J�ܰ��!���i�r[m}wxBǇ�i}��u<�>�X����XӠK��Δ�n��I��O�^����_��vv�����\�}�ņÁ��a>����{��&Ӗvm�����.�K>�N@Vz� �O��n~�X`��X8X�T"K� �/�E�NW9�KVF�t������GH	dk�t�V	U�Krr^�i(8Ex �(��z���]Z��/�∏���zN�V1J�rr�x��7�h�D$W���ō�E=�lCk�&�$���
\5�w�U�PX4��l��ֵ�ˍ"(B@N�h�t%- c�����A��x~䰞�x���Y���W�%��E�!/��<v��gP���E)��5,��w��\���H�A��J����J�s��_��Y�u�O�YZ��h[�V�_����P���( #�R/̽�!�܉�4��9��4��TPm!�?k[���$��8*�i�C��B����T�}�������{!�'�%�!��=\t5Q���n���������CdAf�5�׻�gk��<T�Qi�T�w������ygF����Σ,�)
r�o�Y�BԢ�e4H�Z��TZ��.�7�w٨J"���W�^�7��ϒ�������0ѓ�Ϩ?���z}xH����߻,�6e���i9�Pwҥ���㈒���z���b��]��%�G/���!7b��/֮�ҍ��EhE3�~���
�qf���E��TZ�q{�a!���j���X���r|r�\�C&�����w.$����n*1z��4�4�������%�2m�=x]R멣�D�9�C�$�b�A /t�)f>ְ��d_��K�(#-+�^� �����-i�c=]��J�
�P)�5���Z���$��/h��koA5��Uj r�\t�3�$YM��Ɲ�	�)c/,Y��^�h0P:���!�%̙��5�Ђm.L�8��M�0mXB6(��Gg4�5A)��N�u���B���|������9]+t���㥯���ak��V�Q��1p��r��]�X)T���CbEI��W�r�>�\�$|��#?�J)%������b!9l�k��&R��Ԇ�V��E^�����r��3'��X)U��ζ�pVKx߼#"O
�9"ņ��Y״&\������<K�����vr��-I�y�o@i3�*?����8�Ϸ�?,s|�H�FM�j햆X���i��ӗ_~)�ݻwO~wvv6G�|��&ʓ��3Zͦ�z��%}��o�g�}N�MF�ޘ�<����+��7���z��PZ��@�(���e1�>�O�?b7┾��3zwvF�����v�H�c�Y���LbH�5}G߿:���.�ds��t�V��;��P�5��+�'j��@���\���m����%-�Q*�
i��b�е��o� 6z����Ƀ:�����	�S��#��8@�$�͓�C�0�X�{�1/NgzL���h�қ��k�,��ּ2�fA�U6�5.~�Y �
%��U�X���Z)�qJ�0rm�녝�I��qyG��P5k�:�<��X�O����]����Bv� 'U��#�.\c!��B8���'��%��*!W�H煰���kުT���HȖ�ؖ@mZyM˰\䵅X�D_�$T քR�e(�F/\�]�E�h�g���E}8K��Ĺ��x��.;l$a��E*	aQ�yAu�Y������+��F�-�\b�����"�]Yh�,��IT~�c[RM_�s�x�{��AHXNC�7R��B:�J�bN�KyO�
ׅ���̳��{U����3G���>LX�]�qUO��D?����������?Y��BKQ���VA��T�6
K�A�S&��g�6۷Y�y�:s=p��=�
���g��:�����0�/NOd���ߤ�ϟ4���%�S:}H��Y�;�S���`ը�<1�ص���(l��[�l�~����_��z��ys�����ۑK���mE��¡��?����t��Mz���%#>~(��@cڻ�K{�ˎ`���N2yX��hp��� K
�S��݅Žea�٠�ނ�Q"�����j�-�>���y/	7�r���vv�E�@��<�7b��J���(%P���t��gl��/Wt���Õk�d�!m-~=UV�BP4�X$���Ե�*��F����d���Jh�EE����:|�XR������
�jH@\����ܑ~�L� �"
�ņjQ	���"�3G-�j��5-���m�a�v�[����ۨl%7Y�aެ^l�� 9�ŗ�cQz����/�%�M�Nщ��s�,o��1�G�o]�{l[��9�;��b���f�7+q`�s��ְ�YmЭi%���k����J)�R��b.�p����F�u��R�1³�y���q4��fx��<�p
*�E0��)�����<?jo� ��������N07��f8·M���r�=6�}�򳢍��{�}�s�{t�x�� �����ߙg�Ew/�+�ϖ?�����ӧ7�.p�l1Y���#�}��C�.��+�%���-�E��N�N��L�O�[Ѝ[�4���Vtbh�N�.sz�.������6�s��=B0`�?Hmw��-�s��hA����z�?���1��(�ݝ�$c��C�CcV��{��B���pE]ibB4�+bm��8�邿��rq���L������=�{*�<��ٜ�Vit�e��#�{8,�7���.�M�r��kx��B� �<�
C�}κi&�O��V	%����R	����O�XJ��Hf*������9�Od���E��\�/ 5�_R�a�kx��o�ED])�"Qz�vԢ�]��<�,��z�K��pU���2�޶�ĺ�Wkmy]��l�Q����۪Ħ�"�ݎ�ӇF�7W�����w)jV]�m�^�=Xۜ=����|���x�A�O_��\,�1i���-�υ�M�]w�z}�W�6��A+�ކP69^l�h[ւ�����T����m�Ȍ1��������˞�F+���s�B�j^�T�fO`�lQ�u��mG,�N���1��_��N�NNԠD�(���lA343��8�`Yu�E�c]ܹ��B�����	@��S�oR��>>>�[��,�ΐ;7YF����TQ�<�aW#���#�ycB}>91�$�P����ҷ��I����'�ZLi�D��v�Z�
A����N����r	����`��Pt&�q6A��E�v��v��>����Y����{t�B�ۋ�0���
��働�#ؽM��V�)g=M
���yO.��f{���B��6l�_�^�nFc��=&��\�9�Pg�Z�R��و��"���u��sM�dZ:��+h�v	�#sF��e�[aY��u�؝�)B�%�4|���ΰ�����΂;f�=��^�̐��@�F�n�Bۼ ���Э��Qm�:����WJ��v7Շ�x�5�@�����h�#^p�6�� l�2<V\U^8V=}����Z���U+B�G��*�{�����\�v�ʋ�cT����b����[c� v�y��k��CJ�U���9U
��=�.Q[x�a�vS�N��M��՟�u4���o�i��iq���[)v�wZ@U��W�y=����X�c��=��J�����H`}�|�P6O1���|�k�S�3�o�A�u���١�^���/�����݃���cʮ�t�qL�9�cА�%+�]��򿷧+�(%>�S>�CQ�K#ڡ��%�7+�3�w����\�B�d����Lܭ�W	_�ei`�1��L�Պ�@-�dp�g:�P�*���;��'F�		��x��y�{0XP�n���J��B,Yj�S+���!�{����n���QgM��:��C��e��あ.���y�a)�,Y��14菄��+��Y��(x�)I��N[ɥwŃ���?݌Re�,���5S��Jxŭ5i����Z�ya�g�����	�L\�1��Z�>���T�F����G���8$}��m�p���Uط���wqY!�4��w%�^\/�ʅS[T?$���_OVchl��M�]�U1������oJ�{�B�D�H��v���EC*��*���UW����J'lLɀ	�Zi��J�!|��_�Ei՞��h�{+�x4+J�+Ö���:��-�ָu�BL}���5V�+*�&���0|����5�`� �<��{~u��cO�����"��3Z^��徖F�0 羝d&y�(J��0�\����Ӝ޿_6��{����,�o��Ea���L��g���^�~MX�(r��SZ���:"���=��$�[���&�m��4_\П^��M�,�zt0��������~Ib�3g���&�;���X��Bvi�Nh��غ�%ተ�B�
�]��j�.$ޜ�w�j�k=P�h�,�J�Kʄ�%�d�\�:@B�X�Q�B<4��$�Eo�|2�B�c�!J�Yq
MBQ2��aE�
q ��x1H�mu��|ƸX:�R��u�.P
$�fs�����p��p�=^�u�x�#���Fe���oׄQ�д�}��h�mڹ���<����s���>�VޣRY���ބUχ��|=Q|����}6���`��x������R?�lX��(�z� ȑmN�Ң5>��ʧ�h�B �+C%q���RQ��+�Ur-��� u!}���UlYIY��zL^�J�쟙��Gl�ǖ��x �s�s600�zj�W�͎�!��ҋ+�AP����}��:��0�.�������'a�ί��Uq���~�q]A���O�^Ɠ���V��7=G[6��s���J�D@��m��S�����a���<94��(=|r��}�~���tX�)m����޾~C��2���O�{�����+>�+������tr���|�l�#��˱�^���rJ��@b��O�|#]�"~|)l{�q,���9��h
˖-�U.9T <�����V����+�{-m��`�����WL�ԅ;`�J��@ڕ�p'6�����t�V@'\�B`�$?���`<=��-��`�U����=����~�oh�R�:��c�a���@�|?�����g:b�i�&�����$����hщN._<T+.q�w���.	���
�E]��2p��������J��l��H��ϐ���p�V�R�V�B(�TqJ�p@^���~E�।a@�%�]'��������ÖX�+�Z]l����������e5�a��?���S�ѨfP!m|Ee&J��÷�|�5�U攌
�FR�a��kI�K�D�H��d��﵉�B]E�?Յ���^�|5�����K�M���ZL�[v\���C��sI�Mm6/����*j2�w[�\L�6��C�*�1��A�uJB��K�׋��}�l*S�x��ŗ��>6�-���7���
�'�����t�����	^���O�ӊM��ק����*�s����P
i�'E�y�^�Hm��)x���~J{#
ťx'���R�0�.
TX0NF�ZmX�t$-q�T-t�Y��+q�D��7`�(tS)�fK%܀�����i�o�ܨRCf��K���n�u!�̵.��%�充|B�������=����l�e3��S���H�X�2K��|�S	���E�p�n�8�{@���`��jh��P�)�r��qm�r�*�>Ȍ�b%76x/�k�`K �d#�Dh�{H�x�/��X�ݙB���㾺=��.]]�#T�{w6��os0�h���l�[z��N)���+c�E��%`��\�ס�J�,�nn����B��M=��)k�Vly�uA�p@ߝ����
����W�ܛ��E�.6T���� ��yN�m�
;�MuA�>��nrh�`��yi��y��5:�6v�gP�M�^�[��uc���$8CD��yo΃)�5�?��gjZZ~�'�뫍�
j��&�Iv�H�5O�)	��/���$�:mM>��jb�^�Rs<�o�������e�=?�GDBkE'��=���r�}��!}�Go��Ѝ���l>8�j����9��>�ɧ���C��J�T�U|�tuJ�|З��t0����t^Hu�d�0	����&�������Y�nЉ�̨�P	�C�~���F�V9щ-��l2���AXfw�'D_p1;�P^%��,W<4?Y,6�f��#'�M&�
����/���d%�xV������<�&	g�@� �Z�p�!�#�5O>(�5�r��j%�����Y���3���]~H6զq�,�@�]�t�q�*G��>���B���t�Bo���-W�2��\9��dQ��bV���%��f�cJ�
⛬��y�X稈��'�2�P�j&�t~�l͚�ߕ	E�1�����-כ<����b���Ϙ��#V�Ǥ~^���yi�T�kiQ��Dy��r-oQ�R�Tc'���X�����ZlGZ[=&|���u�-�v�L^M3~5��7e<�������J�q��
�s]9|��
�i>�=g̕}���3n>�n�"L�=��׊�|Sx���J�R��f"�z���Wm�+oP|���t�*���V	�����KI?搅�Ǐ���o%3���)�8�G��4=�dAg������3�KJW[:?��і���4 L��b���AL'Ӕ�)��-~���>ga���N ��I��4�*�0���4>'��X`u�t�ޠ����"������+�F�&+A:�`$NP��&�^���|?+��Ar�����L{�n7��]��_Α%:}T�%�+(L1�I�Q�YH�9("0;"����f����F�4�@�5Ie��d2���\s	3��Q�����<��p�+����!*��8��%
�&Ilu弲H��oc���,�#Zo�ReA_�9!�0LY�^�I*Ю����F5T�We-��J^�����@W�^W,&�*� ����Gn�
N%��K� �
��|�V�2�ޅK�@�y��"Jӵ������Q%#ޑ\�*+=��hʿ��%M�ͮ|/}Dk�����
���u�`�yN��/b�-�)r������Rl��kq�k�ۆ,�{7�Pa��wղW�^�}��ź����_�YM�9�z.��:��uB�*𠩼����L������<*اGBC���_k��p��أ��?ea��^��Ź0����ӳ3���ӽY�����o�2�ݼM��S!�8��l���A��,DQ 4]
����t�B��H%�{�$������(��@8�U8�äT
�&;���~$EN���V�I!���07~9K��p0��hWBE���Y��a�VHAY}�o*t)KRMD��	�w�qyb>
��&�n��
w�>Q�<[�g*wk�!��]��v�ޛuިԉxﱶa��;�9���KA［�
��ޝ�{����s����]V�=�vN[bE���"Py�2�i<z���ѯ���X�@��j�3�&ͦu6J=�5�nm!H85�+��bڶ�D$�[�y��w�����E�LI��ږ�kV�a��BuR9"e����TB��L��.&�WO����w��T�7��7��s�{ȧf���q�̽��y�w��0%���U��㄰G�����[�zn�[jX��	���V�.���s��V�B���S�yV�F�yx֒�jT�%�q[�������Ԉ�Wk'��gS����=diy��y[n}a�_���G��٣��_�?�������~Aw����Rp�xH��Zn~���鳏~zrĿy'��6��l`[�k��[����w5"�b���tN�@��H�-R�;	���)K���fs�J���Rց���O�<��̖Mh����V;�@������p4a>����J��h�#Ԡ���J	*�ȭ4%Ggtb#���&F��h��'Î63I]�4L���-�R<)h�̷	�7#���(�B�����$u�pǋ~B��N�\;]E�^/��g���F�KZ�3�d��7�oh͚K�W�b�Z��؈�����ę:������IXs��+��	~��+1M}�X@��W^�s���������'�E�@��6��Z5�Z^_[�/�xl��q���6N���g��C�ue��TŹSJ�SF�7�]�,W���i#��Bb?�^���Lq�Qv9FVy����+	_��W��T)����(�O�k��$�T�&(=��A�Ug���J�CG�����|�.r|�m#�'��y�H+�}��ֺ��[��P�Gx!\Y�Uet�����$���k�ө�i
(?�8��,��U�����qa��0/��I��������W�#����Go���紷�+���E���!�\� ;�u�޿;��|N��L�'Q̂r0�)��PV��v&BG���%�^��s� �:�	��lߨՆ���	�h�-Kc'��i(s������MC{K��Xl`��/�o�߯�/Y�n����m�����6UK=MK%+ ���ā������ހ�����],��8R�@��3ш� �����R��H,���kifD��ђn��%��b��:��ֺ���x��E̸��5�բ�Ig7���Q�3�U+�b���&��s��%	�B�W�z�d�
�h|	W��T-F!'������W�1j��~q�7�M�R�Pi�A6�ek?�*35��H9��G�k:#=�yg���yy�Z�K0&�nSV,oF�Rc�j������>R��h^(TO~�h�l��:����s�o��k�s��"����P��2�`���;a�_6��O�g�?�nHE^
C!�W�!�C*ت��'"�d�<��O�u�ߏ�KJ���hB����d�u�xm��ʭq=�pk�ڸv�9�� �Ga�BҺ��J�a��D�|�clYv�P��$��g����]�]�I�XگSW�\6����6Sn����l�1��)�$�>������r�%X�乸r�3���0G�=ЂY�5۬�<�j��x7C6��z��Q�Z���ϟ=�O?�_����W���B�>z@�~�	��.i���7�a����SIv��y��L���҆�B��,.W[Y��
��#��[����N�4 ��.A:�0aA�y|Vi���O:x�h9��f�'le/�{ĆS��Μ�<�D>�j;���'^.h�Q�)�������[�ީ(�`h��B�+�X�(����|�ŵ�D	H˺��S9b���3 �����(�ۻRZ�ȿ'}�I'�W�jk�����1.| R�Wr���v�%e6����Xک����<{�q�Q�^EBgk��:/���;A��l��z"�XMR����'Yߠ���C�N"���l.RԂ<=�x����^l%|�T5~bC��J�E�WVd�
d��
�*DZʊ-���e(Qі���́�*�����7R0y�V���,"v˻�E`Y��y�����y��L��I5D$�I(� ����N�
����V����ୀ�@�b����n��^aP��Hdg�[)$�$�Jx�Ŗ���u�1.��Bw���zE���7���Ƒ���$��/�2���
�PY8ָ�Ľ��2H��L����L��H_K$tr��%i��³ci��Ґ/ �+Η�)�.�Ə�%�3u��(����MG����jJ<>V�C�$U���͊�Hd����p �6᧬9���D�.%��e�$hl~��4Ixd��/[&���6��DE.��P�o;�;�T��ݫ0�m��U�ۆ|�a���Prv�M6� ���`0�1�-���u։�,���	G���C>1��1y�2�� z��7��?���n��{�o���޽z��^���>�����섦k�rs���͆�O��0�I��{J��^+�|�pF!�;DK!ݓ�Q�s!G�o@�X�dX������~Qy쨺�h(�P͢ �+j�ZM<ʣ���x ,��\��"H; ?�i=�P���:����uV����/f�@��R��-G�
a�L�L��xV�Tm��;���u]���
�j�M�29'r��E�f.��x�R-R�.�^a����	d���gDF��(<�r�� R^�J���uuV��&�$�H��K��I]Bk�M
0+^h�� �����dc0c#*�����Z0�1}<�aP�FV���ڙ	%�g���Q"�`�X�L�7����:u$���Sl��י���LZ��)���� �k���#�U����4��I����Re�v��ıq�,Ԋ�_/���L��-�9���M�\�J�9/&�i��1�U豛����+Z��[��{M�q���a��o�������8
��А�fU]O�A��X�n�(�dY�a���!>���V���:��k���/L����bnM�^#G0�@���r	�m�|�a1
��2���5�g����c��m���?�i:�lsQ���x�������ϡE�:�W�׿�r^�c�}��j��3.�$dgA��Eۑx�X^Il���<}�&o<�xN]Q�Y��z2n^�̅����((|���&ȰZacux*n�ݺ��(w������,Px��ݢlӴ���y��Ϸx.��n��'���<��i�J���5���xLx��G1�ǈ�����B��B�O,������nݺC,�;�T�	i��ONN�ك'b�����N߿�)�$���N�B��>����ә��^,�!p����HabSVlU4�^#�V���\A���O�W��O��⺥.mm�iSfr\0VW�.�lу�5�@�:��x�Ufƕ�#��� _[���I�gXY�P�rW���C|�6ݲ��f"���p52,��FLq��î��Wq�bS�B��$��қda��"�An,A7�I���0B1޳��U�E	rKh��aF�IPN�2+�i���d�ϳ Ȗ|�!���,<RL�A�tl����0�De�yC����/I�%r������7U����7���3��ͷS�ߌ����K����^��7���>�ϯ��?����d���?���Y�v��������.���/�( p����Ѓ�[�����j_�˯����*qg�}�U�t�k����5B���i�����O�����T�EY"N�V��MH�f$:�!m�+QYbi8��rX����$�lE�>H⊑6Ԧ�9B!V*P3WCb\���n��PQ�b�I�F{�jB�J��|�H!x҅R�4A�s��IⲪ ��La*~���H�/1KV�ٜO�.�Э]C���	+i6��4���^�L�����έE��H�K�W8�yjѐ˗�`���HA��ɷ��d<m�X3�;cH ~��P"1�������X�鰺f�|h���"�q�q�q���~�ߤ�M���}�?�����o�^�����P4��'����G������Kzwi�?�{��J�2a���Gh�'��`�7�B[���≑���f�7	��5%,���
��4�>��a!!X-`��UQ��A^�N�d�B�P"�@�x�	(~E!��d��:A�]��H�oy6�iPi�� Oqi{Ο�|=g�
a�`C>���� O*T:�!B��MW���@UBO����>�B�|��-�����������h=�����@�'�����G���C:ywL/�}Aw?��l����#Z̦t~�^�{�#:BW�H���-��kK�)��s�!���KL�<I����f�P���?���b�h%�b+�y�IQ8�[�m����m���.�-HN!�����Uf�S�ܿ���ؘbʖ�ֆEZZ��g}1C�!ūa�7�h�tC�P�V2Z�n`}�U�sE����������l��_
��P@    IEND�B`�PK   T��ZN�v4	� m� /   images/91e5cd07-2a88-4b0d-9128-72e2f992e16c.png�{eT]�����ˠ��Kp	 �Cpw$�%H ��'��Kpwܝ�y��_{���9s���vUݺ%OU߉��*��F�  0d4  j  � ��B:��Bt�R��`�H�oT=w �P����S�^�����t���6s�X�Y�Z�[8;�譅�(ʼ��u�����.q6�n5&��h��H��tҠ��_���o_���ݰj�9�j`@LT_�Z��d���BX��%����T�^�O?�ڻ������;�^�t��#{{Thm�+��j���J;�?��G,d���)���'eH8����%cG��q,%5'��O�N-J��dj, 4��v8?Y#�0Ӎ��?�`.�V��z1�O�������{W�8�^����ap4/~b^���P��^���}��@��-:P��:{1��ΑW LQQ���Z?���U>�Z���N�1C�]ɅS7�HM�3���?�Y0��sZ�ۅ'� ���%,҄nl!���wD���`G�b+��O�~������)����,�J��z Rɻ$�-�TR�*Q8=g��?�Ѵ�Y iEH$#'Iz�oY����+�a8=��b0ҟ�B�T��}��;5ʻ�;$"�;W�P��$⛩�4�_g�,�� (7?�Ɣx0@b��awr��`��1hdb�Ծr����Cq�Ӿή*�Ä�݋�q����LR��\�v�Bo�`�z�̐��I,���F�4�!�����!�
@�p3O�ij���0.����ZeE"�X�%<|)�ؤ!�`3�2����a�ƈH?��¸�$�� ؈�H�QGjC�T�ژ�B�`̄y�#����vm&��"��[B��IL����g"����RhY-��C	�
�I�H�VAt2�w
�Z5����얜����e���!V�?���>4���>*$��H՚�n�	�RBx3N�K�#�u��_�u�a$����8�d D��1�J3 7I�*E�ưdB�������ʠ�DJ�~7�S���yj�d,�8#V��K����������,�cʪ�c��C�������b��Z�8]| d���f���g���sj�=�� ��x��!�&1�r�Ӕ�`�co����#��&�Q2G	��~��^klQ�0>�s�5d g�B=�d�H?�JsVP���/�ama��&��?X5]�(b�Y���ӣ@��w���'�.�7igi੅�)0��VK��E�i*W]�Tu;=�,����?��7q.N�;�.��ڴ�[P�B�6��[T����*.E��ہ-��'_sI4�Ҡ����:���=8R���	*�+��t�}�k���7b����{��>҉"�T>CG����WV�Z�����Qʈ��^�	�?��9�̫P/H�"��w�Z�S�;WT�x�6��:��I�R��E���� W�}�}�{�*К�ì{6\m��%k5'u�A�lK������l�	u��4�x�J�r��
e"
��ו�+)�3�+�֔�OhԠЏǻ��qF
.�^�TȦ<�dJj�_y�8=r�v��g�E���0�ۆSkJY���{��u_�#��H
߾��92��8���� R�b~�4u1p�iF����".pP��j���{�<���ٿ��Pu��,���t�ڰ)կ����ݵ̷��xv�լ)���;f��h�N�y��?���=E,��&&���;�"j2y�0R�H���)d�����m ؉����3�.� �U���ցm�l'�2y�1����&T�70vႝU_�X*�X��ˁܟ룽�����<׋y(a�Bᇇ��|�է�/�Vē�'�)�o��@i�_Gx�����I�UeO�Tl��	j��#��Q�TӃkw���G�C�#�X�ƛ9����2 j����J�xQ�eC� H�X�f����t��tPԯw�A�n�r�7}���R��uNOǈŜ.�{����U��	��z��잤�a;��ب	��2;�<�U���[�0�6CZ�zP ��$�;�k���1�����-��&}��ܢ�}2Bsh�쫠R㥭=�?��65$꧲
�Ɏ"|��b��{����|���M��^�$�0 q�$"��Yo�Mp�+�ڊ2�#⫩�+�>�����J��t+��)�W<!��K<^�>�ې���YO=����Q�%�rpb�Q\G�vË}il�
;͕`N����Ml���`Q�昷�;��O�S̯��O��R�>�}�Jwɑ��mq^���Z��o
~p�EI�DŢ7��M�������SI��C�2�YWT�N�I���#��
O�1 H4��\ԶP��@�^bG�A6~/h�N�K��'����"��Uo3�0��i�ZI9V~�9�(�<�Yk!fӁ�4B��e���%�jכ'>�4��?Hĉؓ��8�tˣw|�AbH*:�I��-FѴ�����M��.�����`�(S>��H���ϳ�� 3�m�j�=�r��.��fm9�B���!�+�nc�x��#�*����k�S�B�������ug�.U��?_�}$J���wB�`\��PL%���17���/���[�YS>n� 0^C2 hs��Vw���/l|���!��}#Vs�s�㐻W25��G���c��޷Y���LU��P�&�:����-|ԩX�z�Z��WM;W���*l��@;���Mc���x-s�������k�*��}��Y`}��� Mx3B�CU��_�:������N�%��WO^��b�*�z�oə�h�B�cNE��<���½׷N_�}�������ڑ�)^���L27oL��Bj�q��Ǒ�9��=(�}���s���=��D��	.<G����ׅ�!�8��t�v;ń2��Dc{C�-Q�g&#SN���Ō��_ -M
�㘑8]U����N�˳6���/E�`�G��f�eG�q���0C���g��2��JY�!>r�D�]
���~Ӷ�$x�H��C$c�pG%�]��� ��,��q���=5�f)a���1h*k^��G� >�s�bQ�E^��J����1�uYL�:�
���'��s�!�9q?j6\(�x}��c��"_�[C?i<=���)�v�e�Uhy�Q~�g��
]������F+9F�8�FƐ,�D��觬�B�.�1	�?O�y(�D��y�Y��"�P\��<�[s����c�U��ߙ�*Z?�H3R�C*Q�����-ȁ���*7�HN���^gA�또�s�����`U�D�mɩ�V�-����i
z�8G0�U�d��;�H���X�95��YE�*�y�Ħd�{|ej2}�� ��Nd��tw�"t�h7���"(�2�c�G��ɩMb�jj�t#a�G�����A&��!�Ԧ'�b�l(��E��4&2;��l�(>T靳�.N �+�F�����U�;��}�mv^�2�vd�Ϋ�%���N~���d��\��U���=�����3��]b^~?++�����3�1���8���
�i����d�H�K��Ѝgb���I �5���ҷ}+.�
&��!�25���Ք&Fa�7�0@�_����}�"Nl+�q���/��&qY���G�5�?(*�5fvD)TP�J�S�Ȉ��PW<R#>Y���W�l����<+V �BE����֜w��]�/؛.��ׂ��{�K�ޤ� EO8[+��Ӽ� �)+��4ro���T��`!��'��%�յ�::� cc�ٙ�M8��g��J�t-���k�ja]�~9:�k�W����t�+��$�]C�3��i�޹��F��=E5�Smi�?�ib�3����<ȯw|�����^�|�^D�7��[�]]j޻K	$Á�P��&(�MT��"�6r%O	�|ԯǳ'
�7-���;_���κ�9ME)zJ��������Zc�T�������7P�Lʀ�DyP	\�Hw2ny��S���J@��E(r�e��Wɾ�����s�R����E��36:duǩ�bĖ�*��~���i���}��;`''œ�§��Ξ���{�5���ɶ�%�Aj��K6��rባ����t��A�x��9��{�i�tCk���D�ٍ���a]��Q��_L3��|�wϥ��[Pp@�G�2
>�ʁE��F>�N�\Tzq�Ҋ� ���#`Ax��<)h��N`\���A�6���ċA���.	��-UȈ������ἐG=-�|xȤ��9�����-�q��[�?�~�!�v�;���;M����O-���Ѐ��3�HM=q�/{!c�� `���|�ү�*OK��0M�t���"*����_,�U/�������/�NM@�n��_g5�7Pi-,3�$�J��z�#r���H�#�'&l�ΰ��D�8U����2i,����V��{#8pB%���eq}�쉻�� k:PJ�Q�C\��𙦟�
���F�=cI��lv&�^��Ɍ��~�Նc���D��m����fWr�P�*�Ƅ�&�L�+��'U��¼�sB_�:`�ɯ	���S>���/Y��cG�vK�O� 8���>|Q~	�頳����p�� �.�k:	z	g �Wq��5r��k���?(�k���R����z�����=�bR3u�%H'v��~����]��'cd��;��֭��G,(y�����U������AVc�m��}�Y!�\�uL��P�b�;�Lyr��Q�"�T:u?��$`���^	�]T���WF�����1�[�����1����l<}<$�i�@2u����`��5��ù�p�\RII #��Xe��i\N���j�X�k?k�R���]���^�pa�x63 ��IYd��HI��&��!vy�o��֩����,�]1���K�}�������8����J���7����j�������u���+��u�$v	���F�eo����J��G+�9\��c��_*q��>����w
��S]f���٪|���(h8Q�D^�:������E�'�e �?�7�e	Pn���I*6�|s�W%�B4s����E<���Ĩp�S�w)��:��@5��솢���YPH2U$�&hh��;���k!tv|c���+�s�h�u��"�]+g��w�TQp��̔�=��k6�>ǡ�k,!�+TEWY �%�b�[/̀�������2&ȍX�*uY� �z-��K�h)6/Q��1���)��Kbldӡ6˟�@ַ��� /�IHۺP�gO��,���|���M�LQ;��7��� ��ޙ�-�x���o����V(Y���ܿ���S�)���i�D��}lY��*6���괷�Ľr���x����.��2S�]k<����G!�u:������AD�8S:"�Y��||�'��O���,$�Z�6C	��X�HD��)}!Hvʉ�5�@C�p��p{b�ň�H|�
��B�}AlJS»k/���^���_��#��}G]�&�6uN+�o~^��0��mQ���G%��[�ö�����r�~��C5�������ͪu��ֻ��%Ց�:�����J��UD}�06��=�[���EjɊ7O�]�F���?��u�-ř��k�V����s���I�<x)q�`"��{J����a.|%=:Ol34��+T
��zK��sN��<���2��g3��6�a��м��� �T�/��s���:}o�G�AE�cQ����o��i��i�`#���\�&W�=�h�/.��قIR@�Z���<�m�ݢ }����15�\�h&fk]�A�ۧ~'�ڑ�CKn[����H�x���� �Q�|�����S$�%�M���bgu~/�@*�3�&�rQZ���HL}�G.,>�g���栊LB�'%e�ԡ`+���X{�(�N�9"��U�~�3�W��?v���"wYz�dρ��w�BJ�̅_�&�7����k��pxMnй�9te^+����@��e��ȕ�o��M��\x|�iW�A�S�'���N-�B#Iq�+K���oY��WeL��OMD��\�<?�nu�>�)��y,�Τa�>w�t
:q��� ���6����!)���c���Q+�u%��p�-��̀��{��#]�p�iI���Ϋ�cR��b�6��ѩ��!��b���O+�b^��|ޭ�PP����*�B|�b��H�{>��}�S��.�Ć�^>O���m��`G1a��HĬy[�LAL�:��V��u% me��P��Tw)%AF�(,��`M 1��^�>�D���-ə��,]���ȩP�Y7���u���C�6�9��4B���>IƐE�v�;'H��2�.��+����j^���;cZ]�Łb�c�;�"��UT��G9������ij.T5�����'����j��k�98bu��o�"���ۮ��RLb@����Qv���,�$pCJ};x7�	6SN%�=�jw����$Z�h�t+��S�̇B/u�B�R�9��2��W9�t�t�.�TJx����)�6^�Q�;Z�i�%��͗e�m��1D��ߧ���ı���y	����#��px[I �� y������)$��4��8��-q�5�=fHz�z@�� �z;����#�ȫ�����jNF��K�I��7�)S�K�V��#���?�?�[����R>����g��9# g�'�~��_jZ;�V@1h�I7�?X��֧��H�Sr کh���*��"�Gb��\T
B���Pq����gek_��x�9�q���H<�iV^�~�_)�B�E�ANW�A�ːKU(N��Z�ﳂ�L
,�[5���P�Sr��N�Twʇ�[sq��D�λ��Ռ�0�����y^���Þ���4���T��U�h���w����>�{�[�c��W!@j�476�B��m�  �t�w�:�G�@B�&��TVXk�ͥr/��F�jВ�*�꩝>o�^�=PiN�cP�U^$�H��M����y������'8��ى��\k�W)�rw�~��+�(��K(ݸ�[��Ҫ��rYĄ�ԡ�&p��E���?άٝ�55��`�4=���O�hÞ���ϛ����лe?�K����/���M��,h�qB�w��5�oT��e�mq���8���k�j�`����BVU�3��e��e���C4�N8��&��p��+�Nd�Y���1��F�]�b��Q8g`}��lAx=,�AHng;Y>����G�Ga�5a��9jh֞�"���ڌ�bl�Es����rЮ�v�i��ٓ6�f��k�Qk�O҈���J'=�)8��Ԗ�.&n��y��&P�E����mc��]Z���x �~sc4���K�+0�LA�iz��Y��`|<���S^K��48�% �%���k,R�7&s�vx����)X
X��8��0D
�B�§���͈,ݒ��\P�T���R��I�`�U���i[`H"@=����S����}�q�=7�胵Fө�_�bo0kF�2���}u�ΘɁ~�G�B��6+��o�́sA�	.H� �|����"�k���;CRu�'�\��7G���
��#����Z�g~[��J�gyq6h��;�æ>�T}c��#�b��ێ�t��jɜ勷R�}���w��o��%s�`#�_�*J�u�>��us�P<[��#��X݄�Ћ��?��ce�G>vX&|A�1��-�!R��6,Pء��a8U�yY���ܡ�0ֈ�B3Ay��F�F�.ۣ�!����U�`��� 0`�W�Z� R�%ġ���孥8R�r���ͣ���E�����e�[4���؄~۰����/��]��f6�Nh��a���B<S�ݺ��z���w)�ЦgOսQ�!�hkN�ܨ����1�.���h�5���U�w4I-��7w}�(���sz����L�=!���r�Jf�å"xTe+^U�)�c��VcY��\O! �G�G�ZpDYY	��G�>�إD럜]�/���4�Z�\����UQa�i��_�F�B�Ǿ���$~FzXgв:����?�hU�J��#�`��YSk[�Ys���!�o�ꇻ��Џ{@T.)IU �|���g�~/��ij�Z@�iK� ��҅M��X�"M ��$&�o�O�1�8�*�܎��9% 1Fi��5Ź����qҹѻ �I���'��u<لc�- . �K��1I~Ħ.�A��?{�0�e�/��������qv�� H�4���v���Q��YHO�����`!Pe��'��st��^�^����GQ�����L�9Ro.��~�^�T@Ot���qrDـ�[6F&��j_ܜc�����P=l3�.���a���A�]E+�dN��޼�w�*�y��`�t�I"Y�v�W��Hhv��%�Ĳ�������-"�/ߡ{�A�b�%>Lfd�C|^f��]F��V�OB�/�U��,�:{L��k˂���W:@�7:���PÖ9�}�h<��@�6,u���F;M���[鈈d��H���m��Yq3��Ж jȣ�����+����ێ+�p�&�_�M[�(o����@G�=-�d�U�����*�pu����h��XV֦�4E���)���8ڮ���[.I�kdP��J��<�~b���k %x��{���v݅��\�~�(�\���;+�j�ix�;_�8o&���FK��� .3کB<�W�-һ�t� 6o�p1�i��޷�g��>�Fw�<\�>z�Z+G���s�|�|�e��Q�z�����{F�=����0m�B05�<�$���k��t�8����m[�%uY
l�$����J���� �u]B$i4Ch�E�1��]�_эCf�lcs�6�#\��%Ej�b���cQ��he(,�=��	�����1O37Ḻ��Yy|��wмE����V䤑�t��N0�a�J3?�������q8蓻֫��v\;��mE��0�H��?��-X{��
�����b�]@OB�����~���d�QLu�>X�f�����P���J~F��B-6��[��#]߳�1�oRl+|Y�o$�O�4��?
��J��������9�B�$���ʯ��V���F�Cɬh�4Pf�ϵ� ��D8�<�܄E{�;�k�]��e��d�A%`�=No�#ɉ��/6@#_��O]���4���(���F��Z0�Q��[ZwIss�d�O �)Ӿw��}bn1"�{vxwU��ŷ� (A_�i�#�m�������ӣ�ϲ'b���v�Iv�^N�ޘci@rM,�#n&s���6&w{'8a��{�Z*�/tAH%-q�,�h����϶�x���󚹯ߍ����#��=J��}Ύg³%F�zo'rC����U�d|$��V^�N����_��ZJ=��=�KlZ1�]r��?vtXc��OqYh1�e�:n��8�I���\Hi�.�{�9���[�NS<���w��o�ꮎ��Vۼ[3����R�?��\!�[8-bw�D����C���_���;huǼq������ro�C;F5��Ng���V�.|�"�D(\�ߧ�u���� H��y��1r<��Rֆ�]�֞��k�T�s�X�YRgU_ʡje�QX-� �4-#��u0J��+ɮC/(>�G�6a-4h˳F��o猙sՐ��ǒ9u�X'+&]�!��K%��~��},�m��"*�����c�·f*1u�ۭ�oo��}���yT��0"%�T�~�]��
��VTdÞ�(!@��k���1{�<��,��rY�5�=�
�V���l�U��"��E:����H���z绡1�w�N4ܵ��"�f��?���=�7�{6��*��D����VZI<U���i�s�W�3�c�ck���*�6]>�7!E?b�3ސ�d�lV���&x'�Y"�fQo��;W��۝�[<�em�y�&��/ʸ��'q��%���I���6���;������r�d����I3���^K��i^&�ԇ�o(�D�{Q~@e��W�*�	���)���D|����o��uQ�D.
��"��\ԁ��큮��[�1IA
���v�� :���<F�$�I�h���S�(��Y�M��Մ<��F,��\�g��ݒo��T.����w߄�LZ^U��5��c�w�
�DN�E��������A;Đ���>�����s��t��c�]q�>p�!aV�U`a0�b�v,�m:v�ٻ����軱W�������n���|�Z^�^���_�t�/���E��`��N��׎��؞_r��j���v�2?bŠ�D�u�� ѐDV�*a���!m�i���L�H��!�a3��/���ߓ�k�;(`W+ k���K��ETѿyv�����P��`���}+暘7<Ѩye�cS����P��*�$E���Cμ������\��ߙX��K+�*�0ȅ0C�s�V���'����J)f������4�՝~& J�جcILZ����6ɲ��H�Z�qD��4[�,�����Q:�iN�z�A�n�=�3e��4����m���?b=8�P�w���=Zl�E��$�ܮ��=��y=.5�/���6��b�J��#?ʀjN��ϳ�?���ęт3����ƨ��c�Ҳ��dL���HĜ��l�9Gۙs+*�8��a8Z��\8}�)�o�&`�r�R�	?n2�dWR�{�|Ya�Gr)|�Y>u��^��+YK�b,-���i�gRj<�{����]8���#�~�=� -��V�T�����8=3̴�.;��U:�;;�n�ii7%���Cд6�xʶ���m]���%T�]�����������b��":O�JV~/�^����=qЂн��	�Ш��olii;%�o�VVb��O���}n����=�Hcy��24ifap��B<���y��m��5/���v�5E�Egݾ�~��Ǔ���Ӣf�����{�&�Iz��N!T���0�|�${�Ϧ�w�`tŹ�pB�����4n�5��W�
C.2��r �s��Ɇ`0�JW�:rajo��E"���ÃR��B���=G���'Ku�ʋP�!s쳚8�J�P��>����Z{4�?6�[�{8V�����P�FVRTt�������y���5�ʲ�^1&HĞ���E}�-I�;,��A�S�%�P��U��v������M����d�D����%�	��k_�:{��TAoz�;�j�2 �����NB�w�O��lx2�Gd��1���b�A���H���]<Rw�>��#%|�����&O��D��|!f�ц���&gٸ扄f~�_�K�j������6Zy���:����̝Ij3�M�ojz|��b��6�P
�5c���a�}:�ڣ&��=qdiS��Ew'?�߅�>|�g"ͺ��n�Đ����U�� �ꚴk	�y���.]�^ň�������k��5t���(�ѝ2��4G�]�8xBa��2�7����<_Z|���ҍ1�;��u�n���}k��rU?�\�r�����ҍ�8<�/���7�7Z�M�G�$_3E�����N� A������hu���u�Z�K��̥fb�F�Qe��lk7�Y�7�[+!��u8����,�Wi�
i�h���Y~B�ţZ�F���N��@�}�/�o�րN-��aG��)��.ua���mRwҿ_��ϊSURrV�^�G�o�AB��~.���,J��vtk�ɛ�Ƿ�ht�ݦ�����ꕃ�c��6�H�M���\L ~�C�b����_C'C}ɤ:�W��TۺW�8�����A=k���#\��d�O�+9P��}�����?�{��D  I�iO0-�n/aX��׶~]>u�keo�H��B} ��ͳ4�Z��l��)@�5��.���I�M����
^,�q(��Bc���?�);�cOkQ1��x7��8W	5��/�&҅l�9|��:��?j�Ǧ[TpW"x��/}v��w)�����9��������썿Ͱ��qp�h���)!�="/ap�.5��GL��(�V�ty�O�{&�)J!ֆ��7=Y�V̧���MH���:��|A��0�+�vq�pM{O����Q�w��t	�]kr,��6�C��3c�ɑ˷�l=9e�㟔�}u�A��R�ѦZ�ˈ�[�_�#Օ��u��xw(�\,=::��m�h���)!qk<"�ی�/��.;�O�2ȏ���Y_�~U��~�}�ҹ j>�K��&�v���X�1�����w������g��J���������67�-�k��$)!y!c�?��7����9
�����]�����C�	j�����{
R/��]}�
�Y���K�^Y�y�5!��R)��A�*�����P�CH���g�T�,�&c��{t0L/D�r�(����<$Ѱ\���.��i���Ɋ��&!�8\��+�J��]9�˔�M "�=�a+����ԗ�u�h�I������8J~�����i3V���ÀM�F��S��FuA�L�x06Q����p	r�J�-�����Q0�%ay]��U`�?~arxPV��'V>َ��,p2FI$�y��dt]�T҂�	���7��� �!��P?Y�~Hs�	�.�{�ﰊ�wy��?#��3��Kc��|s#��#�����N~{.9���
.�H5X�|�f������ ���j0�#"�O������ó��vo_�q��p!�EB���ߓ�**j^�Pi+�Rffx1��%���I����n^#��}˝��O��"���!HܧI��r"��_����W���Q!�PRS�SW�Exxۯ�6�P���|�2��*�V�8ސ��-?�|_̶��o���OC�b�H�Љ�O��ϓ�5K��e#�#��;��!�7Ϫ��h�����zK��k.�&��*��U̾0�d��gƓ�[���%�j�7q��R�����Ó3����L� R?/Vh��kf���jL�Ui��L"�n��~�v!�j���0�.��e�����q��A�U�4@a���{R�E��D�۩���M!'�$�1�9N=����YVZej>��±��3�("�����+�����p~ޱ�r�`a�D6wV�e�D�IN6b�%��+*�������!+�9���n��
��$4pOfkr�n�m�Ld�zQ��$��q.b&�o�Mv���Ѩ��,�^�������q
�r�I��a���i������y�cG�ŏLt��˧���R��*�!b�G���	$�کO�^�u�1��Q��8Zݫ*F�z�Gp5��C����*��W_d�hӪ�F��8<�Ir�p[wf�:o`9�RI��$V��g����<){��i"~(ґ������Z_�����-�l��SH���7��Q&c륲Ȣ�Ai;q���W���{��oqp�T�]	��Ym)%�o�ӿ[�ZO��TB8�9o
C�\��zk^�7����y�@����٥R���/�F��u/��#��NA�N
eٲI�/Y�����d�
��B3�
��'�}7��p�~"Ih�1%.3`+���D� ��]٫���BXF�;�,;�,�����R�/�;��".�6"��ڊ���b�L���?�^66c��|��$o8�ҳ����^8"83�����,����i�o�q؇ڔ��}�|Φ���.�z:�ɽ_A�S��B�+T:�3��E�����8�M�[h�AJ A0�����}5�664��΂���xMZ+�X~���sQP�g�u[�X�=T��aE��_μ@v�I�g��Xi�F��� �#V�����^���ҷRDF7{�z���AF��˕�2-z��au\z��ӽ�6�����=�<�.�}d�fk��)�*�-��;�N��1�9�g��m3:����wHz�mE������!����O��yYu�B��˰�HV�ab'��J���6�T�5<?�Xv�_�(ZY�.x��<N�k��G&IPV?A��2eZ?�*�L��h��5
�V������"��͞3��p�� c.k�{x�l�H[�~���|�GPLY�P/
�H�/����b�!|!��Ps,'UF_I|G��q,�r�Q�.ʕG�UU�7�����`��u��^$U���BP�������K��9��p��1�:a� �j�=�@*e�;�R��˓��5i(���l]e��9B�cqC�$[�vy#7�U:��V�mM�n�D�"�h����#���ez�����	���7{����J�«����N��cG3Z��=���8�ș�����c���Vt��D���3�?�c�qج��-���MS�t�T��~Z��I&����$2L8K��p�7*6:3��:9~�k�X��3�꽹�$\�2�X�����ߐ=������57]��W�S���U��������6C�Aq|?�5�`t{��hF��=���v�dL�!���(��.�gg���J> �[A0ؔs�^�	j�vژ�pBz�[P�_/9-\l�ܲ�X���y�E0��0��.Ż�����~��y�����.�1������,p��8\�w��4Q$�f�U۹{��|��O�)�$�<L�&��q��̔�ԊM��'�!Cd� �w��H/��� -��b�H#�Hd5t$�zi�����Pχg~��w��=����y�vT�<{�35�eR�e~
m�;�Yp3��;m((���;9��~I�ϵiEyWW�%1Y�GU��1����@y+�H�@��CJ	�ȝ�F��3l_ө���EZ!��?����/��9��-�#��l%T�!fJ?v~^D��3��.���+:t�	魩�(�}���zU��p!)-ͯ��2	��] oALЍ��o�S3V�%'"�]�D���H��Y�>5iϝ���F��
�H𡸭�H�^�s�h���1��Z��_4�mN2���7x���@�E��E嬨�Z��� ��0stj���I�1�͖��?$c�|��j�l�	�;�I;%�P#z��gs>�n�D@�<A�h��G�C��q�ᇥ���ux���)*hԈ��춇G@�Nl�b�cԻ��_�a!t"Z)��������O��'rץXW��#]�{ߌ8 @ߠՄ�-�mr�Z<��X�YP��\�U��bBZ#-bFf)\���AQEųmGq�ⶒ*��H��Z;r����� �٣��:���r�b������6(�>��A>1�4Pb�`o�y��\kV�V�G�T�w#���Q��B#P�x.��q�Z�c���-Ex!�l�F��\w���⬩�8h�і�(u�J?���P��OO�F�c�)���r�̩���Ó�Lߥ�G?×L��S|�:��Յ��&�!o��hZ�V�r)����P��H�̙Or���{�
�
��8eq�U��b�?w�����y�vj�%�g���^���}O���]KKD�,�sW�� �ׂ/���z����kok�x��I���SD��iA�<	qmY���֋!��\Q��225t������O��m��"%���)���.rv����Ƅ-��#��ڹt�@9�~X����y�N{��O�Q˒*� ���[hd�Ŋ�|��~V]w~�A�}sϳ�!��ׂKP ��yfb%��\Î�ŝ렆V@[-,j�R����uŧ���C������4��YX [&�����	�=��z�@5l�c1���z�FC�n(�����i����[q>4�ޥ���ċ򿭷��uƺ�tїg�Qt.��\L#��%��U��'�}�G�����;�x��/��ݚ7����M����I�%��jG�&��5�֋���wBQp %"-�at���*���ɳ봭9��8R����y8��CcE'��85�]�����#��=��Wl�ŔY�^���I����`6?�o�lg1�����EEF��z��m�6�C�%�������_��RV�����*-�oo���>�l/z{�5�x�P�7�����o�ɴ~�������c6��＼�F������V�hi��-uh�&��Q�ه;����k���$6mK?�3�-T����� F�PJg���(Ǭ�ލ��yҘ����U?!e~"�cY�Tmv��g��06�����t;�&RN�6C�s�6�Kfj�I�Rs���#ىuh��6��P1
����K]{m��S���,��C�V�rNq#�<�Z����o�n����+����J�^���G����j����,���DObiC� �6�TU!~<2���zd�¥H~<��m�ڀv	�����^���Q,�dc{���|2cy'�������ש�~퐻<9����eqQ�67�i�=,�`5��И\T��V��������L���n�h������W���x9WսY�2���c�<�ϘlB���+�p?ft��6�#�D�����Ű���ҌZ$j�o�@,���ؚ[f��*~��d�a�f�H>b˨'�M}�.r����P7&0bl��l3�y�]����8B��4�1���p�6	�$�<����	���r�rs����~s�вhv�Fd>�������֧֭��}���Q�����6e�@t~`����L(����ؒ��5���bL�n�[{kQ���lf�n��ym�rp�֎f���\;99���(��l^ʞ���;�:��蟇�]J 𵻅^�AҚj��9T���8\�3�����'1Kj��J��	���&]�͂FQW����+�#ke���)��ogV&�B��th��c^!�����+��j� qww����N�����Awww���!����߿��p`�7����U�z�p�.�ۜ��x7%+B����T�K�������+)��(���^����n�b�w+n��=wmw��8}����bY^��!�YbI�o��3�������P� ��V{�Jj�v ל)pJa�nGQ��>��R�d<����,b(K�o����ܮ]	)��٥���.b�~w3��3]o���m��O��=f�WI+*�/���r>���$���"��N�d�"7�;vV�uŗ�z���a�V��=$��P�^B�?��Z�A��>P�Z7�+�Lϙ�8�;{����;�8�$�'`?���Q�_>�)��T�6k|���"S�kF���,<��Ltnĥ��4([C!}$�--�Vsxk��r�%�o;��ۃ��3Վ�i�n�1��&��'P�1�F��L��yfc���-N",.m^%v!�p�$f��F�}���kO7�(�+��YA�������k���S�e������]�Hiii������W..�PT0� ⮩�f�M8��� ���d���8x���)� %ā]�_�~�ӖQ�yv�[�BV��V���	M�-���o�x�D����lxPlu�����@JS��n�DPz�++H_���̙�M|}˫k2�}�D%����)�#�7I"�s'�;NF��)!�'K�IX=�/IB��م�Ӛ���QĂź���T���>p����.��K��( ��=���pmm-���Wc��C'D`l���G[�JT����Lh��7��/?�.|,�W�pF��`_ �D�>o�����0�4��M���#��7��zj�{�޵4%�)tdki�]�>�
���Er�d��:Ҥ�y��[Q[7T=�I��<^H�c���YC��8#�����,������"'�<Pj�B|V�~�Z��؛ӑM����F��x�8b;����P6��ï4v��H�V�y��Pa�---����u	!O��P����5-���I6X����-��yvV��e�!�QN9\�@��i�*Y�!|�QJ-����_���[�X�@T�T�`g�,^F�
,z���%FL�{}�=�W:��{s�l�d�r�a�n��تL<Ƽh�������#��b�����0H?��n]0y��eMt�i����7ڧљ���Ȥ�L~�3D��',�ۡ��n�k
��P���?<�W�6��iI����[Z���pp`�HΤ"�*+������P:[_)�& ����rx��%��￪����o�k��o�uF��PLMM�ă��h��tf+.��!���c�=N_^�ir&�����EH%��B>h�5��I0t�sA�=�u��DB�cB�qm.�/h�oũ�7��K���SsR}�^ę�U�c�Ѳ��А�u����uБ�����7u�V�������0Q bZ or- ����I2r9u5ҥ��sf���ë�����c	
���Y=�/^?4���F��]������F?5���j�U�����'��������tE��1!�K��J=t����M�eԯt��< �ZU�V�:��^$B�sև��L�[��@G�|E�|���/i��}�Η��_���*��JuA8x�T����(nN�/��y�S3\jX$Z ����e��i HD�V��Aa#��K�R���즥T���j�I��cj��sd�y?�&F���IJX_�'v�wU�W<�[rj�,KPLFl�i�a[{��j`H� �0�D+�X��n<�ʽ���"�d��k�O]y9��:���9�ȱ��n�v���T�r��_�x��_�����
�p��t�ܬ�d��<P�OQ�P5ăA5^yՈ�:�!ۇ���j��;p����{T���t���B߱�A��)�s�lo��r��Te�F ���b,h����r��Jħ����zT����:�� t��X��i#���&38�:ː�	�n�Eɐ=lp"�L�� �"��)4��=�����
c� ���A�6��[�1��m�����z�ֽ�{����.w�L���I��k���I5� M��T�������K|>I���d�	o�J���圁�c%C�Kio����y���N�����zF�W��Ӽ �!ˊ���8��<k0���<`����Q��ǖ5鉫R�D]����_!�s��[�8Ȝ/;������	<e���2��N�Jt�:a��V�&��+4��D������S�p�L!�έ�Ǽ�Z�G�Q�q�b^�0<.��2F������8na.�ta}nN9�,rwB���2�)J��5�g��Ks��كU/
Es;�q�k�4",�����%/9��ӗ�&�d�8�b��t��V��ݥ(_���{�K�B������j�,mP3�@��b��- 7KeFFщ��
Z�v�Ŝ��ضJ������!.�3�ʿ�iyԢb`g5� ������J��_�o�$E��L�׼"�[z�OUj�n����߫Ϙ�t"��I����%��;�Y�@u��KG�SOG�1ăVfNKF�SF��Կ�pȍ��Bf��Ahtn%Q��9���D
��R�:��X�]n������`$zm���|g����ؾ�q�K�̄��({��@�iY0F�$
��=�Zi3�qE�,L7���|7z���zј�f���c�znIL��3\F*�Z���9!#Z<n:n��9�9&〪9s��/I0�g.x�NȤx����*0e�b ޺�ĖT8�L��\A�ʈ�(�g0�������FA�Q�a	ѫ	�F���y�e����k<���ۨs����@]��㳻hA��$û��fdk���~���,����+S�R�4�:���M��ú"z02�q<�k�v�ʑ�H���U����p����iLI��Vj7�;���cI�bs7|5�?��*j�\j�ײ�T:�j��\͌L4̇�Q�N\������/��k�`;1�����4 �G�B�g"f����.@AVhͥs���r�=���G�?ت2����S�x"$���h<$��Os|��nQ�{ �x��Kg5�b��D�ڬД��xJׇ�1"M�C�ʬ_��]c�T���`�V\ōy����*B���9+�dqW��KR<�i������r]x4Uw��k��}�FNb��%�qt:6|*��P�{�O�s|�LP,�� FƉQ�La�y�&U-��u���@���Ȅ���p�n^]G��&{VZ02J�%�)(0Qc�:fb�ķ���@�i7V���3�u��q1��\zؾn�Q{\�T��b�Ϣ?P��8�܈#�D����˿�W�����u�tu�S�B�i%D�l����P~�Kt	�iRF� D�1�-):0|� dpa�a��w�U]W,l!�<���
��F�H2��U.��,�r7u���.I�c���,�pV�"G�ee0)0��GA��Da�|����Ad�%����r�dɄ3��p#�#㇀&��
o��1��[^���U
�f���c0�)�L�A�ą�de�(�ŉ5�~�CG�Gxf�Z�#��r�D���ķ�F�S�N��jG>f$S�WF�TP����a�_W4I�*�׻j:�yA������`�j� t�$F�1�Z��ʣ��x�����8M���g�M)e�e�sHR�Jit��cR�� h@����Kz�u%��+���� !�����b >��H��(�`-\D�b0*�(yT��1&������a�����.c��7���v,_4�"�����߽�ĉ0)'d�h��_������H����R���~��=�+��H��T�	��4�~DZ���3�F�����뿘��z��H����{%0�1Za�p�t_OЇr�>g"�[�6�K.�*���+�FNl����q���k(5��F.�豮%�0'��f��Β���&�C����G��p9g�`5̨�gnFR�	��(���;U&}>G����1h�	����tp�b��!2��3�v�x���G��ߡN?�P�-|�ߙhK@;� ��33��<6V<Q�#�_Q	�8QX2�e��%ѝ/V� X>�:�+����o�6h�Nk�=F�YnFt�AKC�i�J����ލ&��Z����rRG�x0��*Ng�ܛk����� <M��P~M@��+�\q0j]�jG\A��=HDv9l����-�m��i;ziZ&GT)�;n.*g۝�ߓ4�ɐ�(���D���	��D��|�E�o�"���C�՜"��)��NF��|�q�|3Q{�(��=�q,X��\�f�s#S���}�MW�	]�:�zO��ޜ�Z�����A4$j�%u��wPh���U�������J?�'�*XPvH�Z�H�̱Mw���L�V�� �&��F��K�*Z�x�j*T�o_ݥ?������cO��
?(т�^6ph���5B�W8"~ȬI�'P�<o��ʱ~3M��)���؃ �1۠|5M #�n�r1��k0B�W(�x]�χJ�Z�͟��p�v0t������� �}��H�Zi�����=H��=>�( �tQ�lCX�W^�����L�d�gb]R%��i���}��O�d��Wa
;����Z&���1/^)��kBD$�N����Iq��gߐ�ˢ:�{�=M����&���%%�����4���9޶M�(8YZ�Zb;�|1�9hfv�G,}���4�<i�ѐ����m~]��M�g�oĕ!^}^e�%Q��$��z�!Ѽ�&G��,��H���F�
K��ϻ�)s��HO_H�3~��c��bj��̛`�]��	Vz|
B�����t%b��詫Q�������ҏZ�b����g6ܒ@�i�=�I<$u��X	��v�R�6��Y��
S����%�O�Jԋ�
��g�/��|��]�/�g\m�I�Rc؟�YJԋ�@��!�؍;�E~���i��L!ar����,��x�o�7�E8r���<6">]��_�BS��&�	6�w����Q��]e�E���Ѩ�E��������� �H��������m1<����ƺ[���Ӥe�g��	�� Z�d���$2
�J���Ot ��NCTj%��,g {P�ɤ�Xs���Y��A��\����Ru �`����˕��/cGI�tE�f�TE��A8:��*Q6�y+�|����P�j�q@�\n7���P�J.v"�k����v�R�p�D�Q&���hMoQ.��fQ9�X�M)rتt$S"�n2��$��եwmSm�Q-)�^G㾌nl��4X l6�ئ�l]=�����rbS*�S���)�#���8���-�x�qkS��~vFj��t��(�fl�v�6�y,�b:���f00�X�,�k�XLţş@<6 KE�&��6E��hOe��z݅�	��̟���<MF���T�V�y��)�%�5$�����u��Q�k�D�	o&�����.=�p ��@��PIϞ
E�i�P�U?�&��2��S�U ��!����<�� O�q �Te�wlᖽ�ܙ�״���>0�u��g=��ns��BP��D�OB��|����<��*�@'��݉f"�A��t���+\�6��뤦LCm]M!ߐ(�35���2,�MT�������VL��?3������S�YI �G�_>�f�76� j�K�� �3�DW�L+a���C�q��,=$����_߻Q�Veqb"��k������n@o<��7e�$f���~�'��I�tN�	$��D���޾没��}r`��&�1tR($q����-*�����0(�G㏃�d�Q?$\���7X5Y���؇��fm!L�8	~�\��9V��Da~f�� L����ig�s����=���x� �84x8R��.�*�O'�OP��_M��HK���^u��x���x���L��X��1ߥϚ��$ܻ��wާ�ʧU�[]�T̎��j�G�u�z
�E��3v���9igeW����5����z=��������n$�X��N��8d�kqOqH�����m%�|,{F�������'�c���[�)n�]�Wm�Z·� FN!-_���X2�|pdCu�ob^��}�RfDy�>j� �JX5�\����*Q�Z��?��"�|��^ �:w�~�~�z�s�|D'Gf<剜i�����z�6�y[����6�"tw��p*�D8����y;E{��~'��ZC��̮Y׍�=C��U��ˢe'닮��ʯ����"��A���$� ��{~D��	Xr�8�L�\`�S�̎�c�؊�Gg��<̊����P� flL�jʹ���*��Oµa��+OȈ��T>=�±S���Ny�:��[��X����~�yC7><��{�h���:�2��26웈�Yk�x�W���l��j���N#v���=bܾ_1��wR���۟�S\k���||L��o��I���v�/���j�{ ����z>�,���D ���e'�v�G\8`k+�(�P��'��h0�W�+̤�j�*�qêSu�h�cu13*�D:�N'Z��!���A��E`���O�5C%���Ꟙ�{�z���Y&���P����?���wF=�o[n��7Y�p5ԓ�U���`��b�_F�U[�`��3ǩ<M��f8��](��c2r@t �0����.N��X_��_�Î�*����Nn��ȇX�ݜ��Y�������&�P�S��u;���s�I�k ,8ks)j���������}� i�~#o�g��~�4��]{=�*�Ki� �!8����=�1b��}�1Sg�2U+P2��L�˿C�5��`vu��� Zv8"T[�r%qW˝�D5L���D'�4�~6�,<T%�\D^^�h��o�1��#)w&�*jl#}%�����rp�XA������O^>�����y��ŤL�e�B���#}����2�=�}<��eḦp����A�Їf?\թC��0���4��3�-zN�o�Xy���rw��e��D�нM�#w����{m���_%�I��%���j5�}��)�9���6abT���vD'�i%A��0��k%}�wT��Ɗ͉���W� ���)dF������4�t��� W�0�=�Jj�\�,-G�Կ�Z	~�2�Q���P�P�iX$̧5�E$�8�b�R��1�7eh\r�+�!g���}�8�429x\˦�x[~�E��I�ؾ�g��8��`�������ha^7bFvqI��;:�0���N�lޱ^�o��?Еh(R��L��ȫ35C�t{�����I��+I�0zu9qII�²�-�e��fh1��H��`֩�d,�����_m��((ŵ�|p��ߙǧ��� ����Vx���[�����	[��b�������+W��ܨba)��A[�^�۸8�Z�"�������Xm��*B}�3Rb���y��z!N�B����%�)ma$��Cp���8g�\��(����'Vk���R	��k��R�y|��#(�$j4�Z�_�N�9)}}�;�+�#;��y(�Z�7`�%~�m�4y�Q�ɳ:K��\(��ݳ��!�H�6�}�ǚ��X`����.�G��1����׻ƒM��	��0!5?Tt$/7�eև2ɋ+jTd&&�y�ާ���5�gw�h{`�݅�\m�l@�T�:����Z�U�HIea���3;�M"����tеƏՌkQ��L�0*��1�6�"+q5H,�	f��ě��:7h��iE��η4;'���\���C`m<���T��%35gx�h�B<�d�P�i�lm�\�y�� KI��Et咿P�"A���l�2�t�����im9�J�`��6�߈y'_ڹS0@�-���7QRhԻP�\^د^�v�f"�>�a$u��-�	�[�[9G=���Z�=a��Ɏ���L�2���C�ZX�G�`�	���@�1���Y�K���S���������t�.���2�8FM��N��g�#�5^.��ِH���S0�*�ϯD��N�H2��ޯ&y����q��z�]%���򢍮�M<�Se����YJ
�;���
���V���g�k�1���_w9o#����߶"�>�/Mt��$�	q��F�|`�W<Y���s�34\��7���6��]���W�Xъ������HH�^�*5��C�ܭ�2���	iB~7m��N�Y�$��E��j��so�P"j܇�K�Z��ԩ���̣�`3gy�ܶK��� �� �ъ�6��g+0���o���t���'> 7�c��Su�����:��CƯ�������_�}V_���Hv�Db�䇪�lu9+�lXN>ZyE"Q�|�$6P��HBl� .���bwN�Xj�'	}���Fo>�]�:�/1qM�Bc�1=AX����l�~��
��N��wu��e�b�ԏ"e�}��n�,�5�� n��b���nwt*�(2���e��/ԅ�
�f��)�i�;�{�60�·��[+��?<6F?���o�~�ɫw2���޵�A�)KA���e��S��_R.#p��6���` �'?Iۦ}�.3�'�;!�"i��_��;�/fq����9E'ey�d�Fr��!�e�S_�D��@�����zW�ER�{>�).)u���u�B�*��w�������[?�����6;ﾛ	�o�����&s��>I��(�M��B��A��~M<D�↦�bq�W$�N�������<�j��M?��,�m����|\��G�OV'ey�[v&�p!$�r8��5�0g�����䣫�����L�P��cl��nv�;���}B��p'h5��C���ˊ@���R�j��O�|4���Z��xL��xx����^�t���.�`3Z��IȦ�.rsRI(
σQ���ri��;����1KfH5�uFEB2�̠w#:4xg����Y|��fJ'�j����&�h�����e�.T���D�.2�x���a�u�%q������fH���D�G��\�'�#�� ���+�+׻���_v-B�Eļ����k�[]v_���9���-��m�*Óf�׳�%��K��Z��ݰoy&�N S�n2g���<R�/4�]['��v:�q#`�?��L�*؎<	����V?hs�4%z{��t���}����eQ����)�;O�>�zbR[O+Ҫi��3=�9z�u?J��d-�AR�W+�,<ؖ����9Ӱ'���Q�Y��9�b��?Y���
��	�'��Đy��Y�v}�X��',b��o�x��p]��	�O��X�ҟQZ-y����<ʵycxU�T(@A�0h)�����0�@yh-[����%D3�V�r���3HP���S��ŷE��#��FtϾ�;!L*,��m&U�i;� +�B<� /��H?�l�`�Y�K����p��8�=���v�Z
�b��mt�&��O��Y���r���]?�1��o�w���l��ؐp����L��V`��d��%餓�&�������T?.$�z�F0C��e�by��p��$���F_�X%ϙ�����������	�?5���ml�z�������xU��~�������ȼ��u����g�����ޥ
�,f����jsU"o}�LGٓ}�^�X�P�x���hM�0�4B �cS1��o�s���ݐ��sd%��Yzl�ģ���9�*`�kj�kNU9<]	�u}��o��B=�+>z�Fr��_l0�v� ,�y]�?�Ѷ�wm��-!쌡Y��[����3��������B���t3�K7���#�� !-ºK!�#8�s�*���Jp�ۗ��dO�a[��[���" ������ǄşC�yQ
��<#������X�����I9-�ܘ+��Ȇ.Wz������D��H�N�7HZDW-QK0�.̊O>ϻ���Pt�Ȑ��B\6z�՘�D|po	�X�'J)Ϭ��1�svTӣV腀~��K���S�NB�83q�zJ�ז��گ�á��r�o�Q���hͧ�|&��0@��S�j���|�{�\'���Y� _9�B�O�P����+���[Ԟ��gš�u��BT}_� �J��A���O�X/��)�p
X��% ݂�	�� �B��
ε�8�s�gF�I"�S�j�w��j�q��?�E�(7kOO�1�m��`m-���K��<=�ѣ�t,��8��?n�zQ�Zʙq�ˌx��A��z���=�E�H� r�[�(t�7��V��K�M_��P��(��ة ��c���x����$L!�D�j/������#��'!킣]�]R0��^9H�*l���ӽ(�F%��'�:��֭�Rf�C�r���4@F�S�_>>��BtU��t�s�Dwe�ި%�������T�!	�d�3sm	���(z�?�G���R����z?X>��0E����6��7����C[�;0��u�����=����Pb2�����1e;> x���p՝��Ƚ1f�q%��p����'ȫ��b'�J��	�>F$/�Fm���P�ˑq�_����HQ�A�i��V.�]�-?�*�r���Q5�����a���c�K v��^��~DS#;�/��(��~�����Ϝ���&e������\��R���݋����^�z����jOvS�F�]h��-a*/��T�J�eFc
N���~/ˑ~�Z%�s1�L��/(R�í���н��Q\���ҝ�u�uT��ܷ P�;1�=|��5�U�L2b��{L��$������!.9���!+(���Z�R�� N�-��S�`�[���^N�;L,8S�\X��s��0�JG#(t��ޜ��ޗ0C��O��$<���\]5u!��i��=)%��L�͹�:��z�t6w(lW�b�Yn{52�L�f�4����
�.�8�ղ;��g �:f�d���r�m�o�V�ݜ�'�	����:���6_�\i
�����b]p�~
 ���;j��,.�������f�S��b�\u��:����Nl}��[��tE��jČ�{/�f8��)b��EA&���@ļT6�axXퟔ6� aRvgjtV�H&�+�K3o;!��Nkz�1����Tk����oN�P����7���uIl�,����̮�i8{z��K�'�U��y�/����,|E7z������zp"�?��z�U���k���|֞wBp�23y��� ɶF�2�(x�N�[�@B��LM�-�K����4!2�����e�h�W����G{پ2�ha\kĎ_T�Mힻ���d�X�7t$�́�__�c�rÚ��P����ƀ7��Yϓ��y�0|�> ��a -�s_��ȭ��b]݂S葩��|81B��C�5����֤:>�K��,GR;>�6/d'�E���(�|�T���^7���{:+����L}�i�.���ʟ̸VF����{�"��v	��_]�z�~K��Z�){ի+Q��'A||���l�/�2�D�9��'H�;��;���`4q������p.���$:V�ʫ.�� ԝ=�pei����i3�m�L���JHAǞ��K~�ֻ� �����,��T4OD�N"ʹ*V���5q��/z2�+�����TO��D����}F
6�I���/������l��p�D�4W�Xѳw�{V0t�|�E3 ��ٺ��]�D�<��g7�I�(V2|�z�[���m���M� FӼ�д\�]�}%5�N��ams����֓��?����r�E���k�#x^�<�5����
ѧ�4�"8��^u�l�����4]H�$.��Y�?�ŌUNT�r�IEq����Y���}�n k�<�����^�W	�w��ED"x��-��ʬ�����K���ZV1oj�0=;�{�����Qz�͚R�c%�ps��VX��5��L�W��L�i��������D�rP�R�3��&��]&|������b�HQML�0#Em�p�zԩ)���Д&m�Ek��B�)V$Sv|7��iҸ԰]i٨�aI���p�D�&0J;��>�P�ɂ?wo`�-��?��|���?O>��R�y���>#���L|�Q�D+���ei���.^$t{��&.S�֛b�;A��`��#YƷc���A\�8���7njp`O��ֻ���9�H�]�O-*ϯ�a�Ajj�#b��������@i�۰R�`�Ǫ�i��˭Xy��
��@D禉c�1C�ޘ�m�+��[� �ǫ���CTw�x?���i�AK�~*��02�3����T�Ԍf͡}��tz]&��ސ �h�n�}�J=8�;-mF& Rc���B�H@<�1�,uGS�O�c�E� �6��Ƌ�tN4��{�.Q``��z�iP�Tfjڮg��JKd�ع���u^.�t;�y2����4��e�A�u\/������3a3a@�I�b��V��Q�2�=�{���������f�>����`��[~s%�[�,�//0���V��~X�8X�v"|�a�*ணf��_��6�	Z�HZdqrO�?�n�-�I�w��6�/u��!�6�j��е�	�J{ �q=-�L�B��t�W��;n#��f�y�rÿ���ĿR�T��v�ۮm��O��=)�R�PN^�������f����z-��nC���B^��0���#����Ķ	e������שW�j�e�uX$�[�s�ß�S'��g� ����<��02e߇_��/��YA�HA���b�
� ��O+=����LȞ��-52`�T,n٭f�_tb$��!���}~�����l�LQ���9y��݆fDp� �]:?��}M���Ǒ`1�^[5���\P�bu��Aч��A,�s��7�#N�7G���52|7��<=}S��i4(�D�K]F�\����9�=���YyT�<~)��ft�>�ּ�,0J��y�Zp���@��.��ΉgS��R���:&��C��+���`���"d��*��d`C�'�]\��}`P`���� ��*NA��hj����E܊���ٓ���@
�nm��J��%s�Au&�%WD��3��Z������BB�{��V|H���i[8z�k�	#���w}��]ZW�b��G:�Bݭ�R%��������JB2֑P��~E���P9������\�d�������E�b��)���g;Wq2���6�=$-5��w+^O��R�%�Oi�^��$ϕF�y����:D?Vi@h�bi��o�P"���t��� �n��=9�{�d6fZ������i�o}cԦZ��~@��\��v�����#�%,��x��Ɵ�����9S�O����`�aV�O�tBw���y��Ƞ(q��"����"O"�?�[�p�p�RF��gC3`f��#��F,O�K%4pp�>��y1�)8��
����+��o���غ���8Ko�8V����}�r �J��L��,>3W��Fd�K�E��Mf�Q�R���١��nt���E�"p:(�-9�Rb�M��h,qU�$F����_����%��"��[ӽ�����4k�ղ��%g4Ӓ�tp�Dj�rs��	�aT��T��'4m1����`�+�48c<?���2��`f4#B��kJwhnw�X�[M�!�fsԃv9�k	�ԂA���EV���[=�:���Aiɨ�TdA�N*b!�~
�:�Zu�H�b@���=dZ�EJJ��YDƀ������ᚷ�s��!�g���[w,�f�D*����qU*E7�cAi�����4�=���������Ax��uw�4 &�^�'�Q��]Niu�ƈd\��NS��ɀfo��*��?Z�T��]�r8�OlW�f��̬�_�ޜ7�fP�c��ҧ|^5�?Z��(ˇe`	Nu}�cp�`A�V���7v�ӑ��yi.r��b�\9n'�AV�j�-�\1�n\���J�"�
e��?�����ÿ��#S�)��kdWb"�c�i1��d܄E����.r06��feܯR��V�ǯ�k�����W֥��L�î�[j`����#˘��HJ�����������=!�'��w��5ր� d��׹����U-�&M��\��=P\_�9zijf�-�{��U���(�Ug�mX�v�s�)���q!u��	�l�p�߳uW�8��� J9��ND{I�=���BhJh%�j�m2{�~\�5(rzӎ���PfG�њ/�W{��/@��0$��q�!��n�͞5���CyƏI�������na֤��P��_N`C����=�U01Ћھٮ���ô
��f$�:��P�k��I��Vg��7���E�dQ0����[)�y�z9�A�v�$�j�w���Ǉ�&r�+#����V�G?����'�B)���OQq:�LBr�E}������`K`��1��z<��HPe#����Պ���Qr��g���8x�x�[�Y�4�d�E�`��.���L�c�����ّQ�d7�jN�CL�	)����e������kM#�^@���J,��K���o0�e����wEy ����}�q�������iI�|��h�������2�(�����6O{-@T3q����7��۷yu#~��j�,`4�Y;�m	�cϷ�v�Bm��8���%��%�A���qo������B�@P����vs�B���h.��@�ˎ3�=`)Ӄ�;x�lk��QɅ�OK��I�/����n^L�����ӵ(�ʝ�b�V�*(6n�q��bb"�W08�ޙ�>n�zj��N62����f0_��A���UE���r��W?��y��v��{&}�`b�Y���b.���,����9p�(� q��~�jdl����o�b��BX�1�OE����Y��v���?��Kٷ��P�b��&(&U=��)u_�_��6h�]���4ႀܾ�U�:$�G{���GYNK�q�j��CP�����X��!�k�_�p��"&�N�*����9�n�#�G nq@=��J+x^�$�<8����SD�x�ޝ��@E���0��e͞�v�ev�<�i��ܫ��|��kb��T���xn���^9�Z�����7󀨟D���d�w�Z���\H�US�4곁�!JbC��[z��^7o�;�{�旞O����}��|�<���3Ç��a�P��fo��a1���c��6ҹ޿#�C�,Ȫp���A���h��.��J'G��)B�S
<\nj�¹��k%j�.s��4��5�}�,Ȝ�B���t�F��"?�0�vW?Nf_I�?��m	:�7aU�z)����thI���\7�޾�T��׋��
?��V7�$�z����ɭ�觊�����
}�S������4P�H��+�o^-w��D�!�Q��V��Pߺ�>@�⺖����s�ϰ�e�g�%��'����=�j�ζg��fďsˉzW Y*��1�>$f Dx��{�q᎘�
s�FKk��a�B�F�aO	�G���n���F��>���0gEx\�;�����]���i�[6ˠK�4��8���;H"���~���MP�%OH����M�Cf��o� ��s6��yq&�j�T歫[��^��A�3�KSS�^׆�HgӨ�4ԃl<���y�Gfmχ�=H���&� ��2j���A�X���z+(��͇<�èb�)x=bth��$R]��# io����m*3I����0�NPz�>=��4D{��3���(g��`���!�Q'G��5�W�_��|��	%Q�#���5�n��D��R㮪�t��-E�W��?�M7�C3> �Bn�
Oy�U\�9�ָ�L�Ń�jm�b��)D��.LT���Ί�=G�A!��'f�#�O^��Ԥ������7zҸ����+Ϻ���r��-�Y�"zk�z}>�5�a��3����뤔F/B8*��!�2�H��u�@�iOd6��Տ��߾�MN9
�+?�etJ��4���;��w�/�J$b|�׏:m�C���MyX+_�鮳�-�B��7w��	�J`��\���uw�Q��(�-߷�ک�+n���G�]Q�� �����
�9Tɑ���YY�^kKѸ!��i������6�'R~�
�Vb~��:��fAD �<z|(�z����T�	-���๦��Q��}L�of���T��fmgm��b���3�G�`8.,�=��ż���쳿� ��rŤS]��D&}>�϶�ܗk�R�k���Ee�{�,���Wv����[�6��U��:��wu.ln̯��-�>f�8���^�ػ9z��pJ��Sz��ݍ� ��	<�.����'�Q�����j�E�J�v&ɥmw�A�ef(0FB!�ڜ������u�m��mz��Dڴ)�3�������~s6(��b�*Zp�,�v�3� 6�``���$`���Da�d�2>z��?K�������dI�e�\!&�vʵ~<���3\Àh��t����)���oO��*⎬nO��z}���$��=�]�z8�OU��)�Nأus�!��
:	�=8���u����)����\��`��<��1��r��4R��Z�{����W ��4�^ �������!������	��w�<��v�|�{�
�����鞖sfzz�	�|w�mw�.��wZ=6�� �ջ��h�<r�x�D<n�͸��^�����\����=C&�vs�rȲ�#�[��߫�X�����u�.X�a}<�h(�/�	+%�q��F�֖1�U����	ފ��!T�\I����.`'D�ڶV�s�3��y��i!*���DL�B�#շy��������1d�M/�$�4�8l�{��&O�f�RR��{�z��wf����'�n��k�����������{j�9їӎZI}�S�˳[M������q5E5K�:�A
��sdwǪ_ie%+�W��0�5�"F*믖��և�H���s����_��-�8ǜ�~��`c+@��7��x������B���Z�8�m���j	�wv�q�!�� ���æY����|�1@dc���$�G��t�B�{PCSPɏw���4�BJ��C��җw��r�Ը>�5F�㺫V^>�G�6lY�l��@M�?D��kえ���>:�/I���Y����pp�K&�����w���0̍[We밚��:𮦗���.Α�\�v�� �TZnY �#�]�&eL����H�A���x�x�y��N[��h'�E��V�Zb���-D����|���x��	���\I:Ǚ3��SC��h]u�%�^3�n�u����#A�Y-G¯�s�����Z݁�����5�ߔ C7���$�~�C��!`�42�o<�!�Dvmr�dXP���y+���:��O��RT�Џ��hh5��x�VeKh!߶�o8Hi�Aꕘ�n��.�qfK��K��^��d]�Jt���`;��AO_9�e7M�4�s�Q@&�׽�L���7^��1J����:����%8^ RS��������{a/������W~����#��6���&M���mY۽|ޓF��I��E8���^�e�e���#x����ߴ]}ᐩ��
��#ף�������N�x���0��C�o���!A�M
�m ���]����>u�?:��zD��q�� ��֯]$
�������������ý/�P#�0֜�l���yno��q�8�GE�E1bE���K�D�5u^؈����9I.����P�D�����A�}:�Q�<~��8��l���k����k��J�if6*�Y3���>H�JZL�#kc�������R�F8�0��$]]]u˧@��i~��=w��x2�̃{�K��wM�9�^m�����.��]�y�/犞"}�̍�v4)�"
��.S5�˔O-�&ժ0ҥ5%o4	��9V�CYhw��KC>�Ee�gc΢5N[}���=q,Z�z`"��h:�
�J�ݽ�ܽ&8���:�`#~>ݎ>RQ^�C�A�ʿ��ڬ���5�o�E���fg^caipL�:�7'�Vwvv
h���n9�ӕ������<�~y��4>az
0S�pRo���(�/)�b����m��I�0�L����5T+H��z�>VĚ�$-��kXdו��!rm�T9bZ�������? �{S����+�l}� �tP��Aj�d$�sa̕�&5Q�3�&鶵��3b��|�죘�jS]�7���9eH�,t_��ٷ�J͛[r�QD�����C�lXp(�w񉉉����;��zY���!?��OQn�A%�
��YY��3���dd'�F�괫eddP}	��f�����Dx�C�l_�޴[��b_�2�@�3+A���YCz�?�X�.k�G�?&Y��`D�؟�L���+nٱ*J]�����q��١B6s�/MT�Q]�I��*D��"|e)��%�#�r�WQ;rC-,[؊j��a�<7wwwS�Y�OxH�E��E�$]D�?�c�>L��V��oʗsF��L���zvnH�W�"r���@���<lדwu��/:�����J�ێ	�q����*�^ ��;�+8��/k�̓�j��Rr�]V�$z?��qD�uB)�<?�d� �^SZ��A	'Dnjl݃�ˋJln+"Ȑ+�4c�P6[*#�kf[�q��j��9ǽ�#�$�N��0�*��vP��x�6AH� 9K�	�ώd��xˀ�'�O��,�Hn�~�p:�9dn)7����5��_�2>i����\�d������<����o�7��9@�y���f�T�<VS�8�By�rP��d��ረ�o�UPQ3��B�a�0���͔+�p�ڎ<��+i��zA�YdA-�-ftH���&�*O���T�˖�7�d��O��GJ]��5wx�ЮI�.}�B��Wuy�^81o7|LT��D��ϼ�l�^'ދK�d�`��X�� ��)cy�,��"f��IL�֥�xgAo+�2Ej����[}K�3����T,���W��T���c届�vc(�	���(�햙MS�K9�廻@���~.2c)�����=K>t�>`�q'�d��O���.C��H*OeZ9�>Am�}�y�{X�"Չ�������uC�廂wN*m�JN8@~��X��bE�$�����a�%�
%[t�0 �(@�ӫ�5�U@7�
T�|z_��/��rY�1	1�kq���}�7����������R������ɘ�t3#���٢���ྍ��MT��:�^�a�:�2��"�ܞWu�7��/�3/;h��a��|9�טL��k�$��ׄ�j�R��G��c�~
v��L�Y�t�p�Ƹ�E�۷<} 9��{-���]�L�A���N�d��++�`g�h���X��#�t쵼��du�.P�� �xb�`�S��H�%;�&H�<,��Tds~G�#D�bF��v��ho�R��}�@m''��'��?<� �#�+X%Xg��r�(?;���ճr���jw�V�²O�q�w�MTE˂?UG�(�"h�.��[�����;�N0!}�J�G�,1/��^AbІ���˿�8���a��e�FY�3���;���܃���J��s\�����v|{����n�(-�1x/��V7�l���
��?��@��}��7�����M]Zk�[I{���x/��KvT_s�	���O�1>S��9�*=Ls��>Ϟ��[�EO���_(�v���#�2q�/��}Eh���Po�N��ozJ�+�(|~?%���'�c���~�g�V�o�9�:���#w���O����-�"��sB�5M�j����G�b��w�`"L����[ȶ]5���.Zs�'F���ԅA"5�zUhuϧ��;ᬿեA�9`�ć	-�Ԇ�l��1���.�5�Րy����삭��������L�B )N�7���Wo.e��^���)'=�h�D�k4��s»�c.h-�����ףc���h�H�l�#
��
�~=���1ӈ�_��-N.�zD�7��It����t�cQ�
 �$!eE���:��B��bcʈ�nM�(n �$
��uZ���l^;`�2�{�wez;`>�����]�F~+��_�*E�r^�xF/���\;lx�N�G7�7���I�ȸ���%�U����C��pe��KC��G��3��?
L6�#=�ʶ!������:bh�?��F�	0?gZ>{ĵ�ckK�g�c]",�l~ $��Y�wl�ԾX<�vh߮��5���dh��0A���MS�L\I���׵?R ��&-9@���3�Ƕ5aXvN3՚P?���~/�2/�]���̟�މ��.ӴQ?�v/���H��/GyԌ�r>��VjZ�%��}&����y���X�-|�x���I~��,��mЕI���g6xHxq�a�<Ȋe��n+������1^[�떵���b[k��a #d�����3ɪ�d��X�+灟�,��]�GO�j���\��/8O:���Ž��l��$�r�_)�:����A��>����>oTOM3�Ŷճ`�Xc^m�Uk0=۽9=[)I���w2��a\�O�C?�Cn##��_��c �U�V��Ύ��E�ыv^͏�F��0hq�}��
q�:>��:��,��L��(�^u�[�P�(B`�GW�"��D�7�v�f8�#$F����h��߶	�
jT+
�i����<;V�t�r��ʵ&��y��+��R�|�3����m�3��k6���L�%�C��������T����3&�}��A �7�N�;�8�hԓ�i�P=K��S���?�4����Lc���'D�V���N=���~��4e[�xV�J	2�܄�`�n� ���e�k�?�?sj��.].^k��tğ�v `A�?N=I*��k"��(�1k�SE��R�B�d��9�\d����@�8	�-��q4��	'<m_|c���Z��|�}�}3\�X������ D�i@��a�W'ǚ�od�����A��ALB31+�Is�(�uׂ���CX����� q�GD�bע!j��G�z�J�|gΞ#�T,���'���u6)�EQ!��VB�Y�ߋĪg�O�KQ:!�X15���(oY��FՓ h>�9���]zy�sSɴ�Y�37� `z	�X�)EX͛^ZLN�\Wt�lV��6�}�/:��c���I�w�����:2nL�èȸi��ʷ6A��%����i��e���Y��_���[�u,�'�M�Qr���V�)Wh0�nk�6���&�׋#ߘX�H��жY|��`hB*��j�RFp����d�Y�Ż�"���'����Hg,�7�-��N%yn�S "ol���{o�F�8b]���j=�N��Մ(���[!��|?p�F����Cl�b��@��NBX��B��=M�.A$@�'Y��ķ#O�(�8F��le��`k@�G�V�:?BR|��.�5>����Ӯ�`�;˲c�&?留8|���n�=�k;�Y�=���`Iаk}ۊ����9x)q���_���$��rP�TU�H�/��RO���~đ�z8	� aӁue�ܡA_�r&�g�J��ܣ����"1
LU<�Sۉ�5��˶��,j� ��8�<��{S����Z��Sκ,(!P��兮��b
�FV���Q#� �
,�W�8������v���(����_�������x����p���Z����"��[e�?,��}����_�9�FM� �2�>�T @�1��a�Ι�=�π���(��@��8��	#��A��P�p�|(�����sA��|��S�� .2��OV�s����P���
�>�P1W]����?Γ���l���U����cX�U�C���J%6L��3���a�f}W���;�&�`:��]�eYX��ri%i��>;m�8��vM�T�����2<�����<�暿���3c����M��H�<��@�&�}�\�ĭI8N�����D>�A��S��PA���I\���6m
s�gO;���z�h?>�KCJ^���\w�L=���\����Q�{��؟f�t�;� ��(���\��~k} �kM��ٸsQЖ������p7�*��9J�y��[������
P���Qf��Q>��ki��R��1�h�d���"Ku4�[�5����G ���Mc��ŋ1^�x�&7��,�DwNFF�y+_Hf�%Ƣ��[��q�j�����V-�Y��;�1'ry�?6�x�����&�Wҩ�"#�Ĝ���
�T�U�Ek��ï�'�������ul�_G������D�0ṕkD7]����_������3�Y#x���Ċ��d_������*���!�X�_���aZ<�8�Y����9&V�9�Kz����VW�O���z�kj��ϿԂ���m$�޺?D,����f�{�uۜh�P�}ݼ�╨N��>�RWjK�n^i�w�YW�H�'�	�\��i��"4���`����N&�e*A��B� 2'%�L���:��_�����s����1)�+�_~�nl5��|D�7�^�E��p�4]W�`EGm���eԑ�{�f��Wt�f?!{��>ߗPi��h��q��fX��v��v��j��e�)�w@��S�O~p��m�b$�+�i�>��%. �@�2Ղ�=���A���v�vK�"��&��Z���$�2�:ؘ�*ĬK-��Q��[7�#N���>���Q.4��q��]��ޢ�!�����Kf�l��p�o��0�,�� �E��v��/��}%�Vޏ�ȃ[Q��_��PUb?�s�g�\���e��.$�?BX�1?�m�|]"�3!�R0�TR��K�iBC�eHX_f_j!�!�J�l`��8���L����Gs���qc�oxQ֬�N��\�y���Nx�j�`��r+p�fj�t��H��$�zPGA�T�8��;���Z�B���}㤬3	K�n�#�ݮ�X�l�MC&��������H	�����}�+q/�Hx���-q���Ce<+�X��2�����n�&Ѣ6G��2�5�ח7k�9��C�ͩ����ɐ��/����*��Yh�۽�o4Kh�"1B���7�LGp?���z?o6���ح�И���q���F�dxm���`3��q�Z�R�:����"����~{Du�[#�P�#2?{�_�*��AnѶMxS�H"�Z�B��C�&�?��S�b5�D���>���WQW�[uLXiC�������<Ն-O	$��/F�՟P|�kA��e
Ҹ�M��]����x橆b�T��C���021:���-�����Ao2jc�
�`bR~`X��+N�N���H|*�@�o�ݜw�:2:�vlV��d��l�k�@=!f�G26I�QX�/Jra�����{6�4QF���^�����G>W"G0zs�qn|�t�C"�/"�1ˁ�`6y��6�����.,��[#�Z��D�����>��5UQ�ذ��-e���l[+S^�|���A\bLπ�P����S�O�5��Rrz�_6's?���jAp~�é���cC��7Y�mCU
�Gd|٬�/~O��ي�D��aˋ����CH����J=������W5�E�f8����n�ѱ������)���ֲ�w��*�A��'qQ�w�����R�x�h��#?�~�7n�����ٺn
4=&(�̓T��O�!NnRh�ciƀ��X��ÃKP�h��Ԃ�Ǆ��"�<A-�DФ���g1���%b�1D��i�����b�[���)~ݸ��	 ��o���R%��اv��?��s�����]dJ���g0�y�/�>�R�&'���c]�+���fx��j�����2�pq��q��%贪}Ra��H�ӿ���S/��[#j1'N���`Ǿ�:<L{8

�>$�����fzW�p�:x����8��\"�Xbo�%E�/�qz)�-[�Gp����6����FeR�ì����Z����'�YK\1��n
�����͜"|���p�p�=˫��~�Xz}Q&�	�m�dx��hL}zq��3{��빞:fPy��h�U��y�ӛ�i��W�!�b<�.{J�Uٜo'��(ة@��)�(�i�i)Χ�z)�zb�3�5��D=1����n��>�/��j�����f����M"Rg����	��Fi���d� � ��L�����SM%�61a���e��]�%=�ɱU����?!��Z_N.P6~=�u��^�o�X�U��%����M�k~�/K��@����r�S�+�����g�v.�z?bQ���q��u�f���b��a�����ݽ��xi�n��Z4�Rmw��.���X��o�ˢ�kM~�_�9+����o;%i�f�Gx���x����*��酢��	b�v�s��k�[���9uگ�v�[���&"��}>�+�?��bV�cE��ψ8��ao�D�szl�V�T�:�k��o-%Ġ�1I��rc�����آ��bKaM�Ye�R\�kM��u9��1+6������p����~ar�b��U3�=�~�䓬�esΝ��{{w����T�Ǧϰ�}EJ�b���'�[Q�σ[ҵ��M�4�l��߶9��	֪6�p�x/.3g� ���_2k߸��o�k;A��P�C;+����KOn���'/���mcN�T���4��t���!'L�L��6�R>�E*w��s%�|�7��[v���{J��_{�XX,����f6]��G��o���Y�m��5i�D��LG�i�&6	`X�	�B.����]��y���)�xz��ܶ־���rͬ�7w�M�'f|�Bz&ȹ�(F��¾�)6������E�ej�J�����g�������;b}a B��:��\���?�ɼK�&XoBj�g���C��]P���H�G����ǁK6U$�\�
	/�����3���a|m��B�Z�]��:����c&&�X�+��NOd澇.t?�u�R�<����j)PH�Tϲ�$��a��t��<��� ˿�d�� $ZM J(*[�
�9H�Ge���@J�M�Fm�X}k��=x��k�����F�'�cg
�1yR
�����"W6qg�� ��a��.�T1s2x�����A;�'��h�C��ɬԴm�*�B� �2C;��ѶL]�Ƿ�!����X��C����d->~G1�F���/�@�����}�Ot�����dj�1:��@�4�X���Չ��{bJR�D=�	��Ʊs�C�+��׵d~���<u@\ө�q:��s�xn�0���^g bs��}�d)�,X�t}����o0�����k1�W��k�[�6��0�V|^����7��2�����l�_�F�]�/0B<Zǜ�S�/ �!��5�`q����o#m��c���-^�j�r��-3<� �����U��88��r����ڱ�m�n���ffOA{�Ԅ���p�>������@p�S�X�T�&�*	�vZ�&&ވ�3y�4<���[f�eW��������&����^����X����d��;ʰ�� ;ݠ���� ��c�����;���rL_�G����6& p��:S�d�_��<��e�MH�~<f6~Q`����f'�ʳ��Cý
����4e��aT�v��*i�p���NB��ޠ��@N����h)�!s5�:�1���*o��i�%���uS��W`ʨՊ������j�G ��sF�I����we�$��d�!�Z4�G �=��HB�+\<�진f�Ob�����y�@\pMr��0ˢ*�#A\�#�^�3�D<�pkY�b����PW|l�=� @e)�~���qG�;��m�'��p��_��ݧ�����gfwd�Ε")��yj/z�l�k�,ܕhň���=�5���C�2m_K"f�ըR�f\��<�C�Lb:u����I�q�������������@'O�/{+�᮸S�Z��F��u
�b���g��� ��r�Yq�[Mr�J�{^��7�h���]���C̬��V+'�ׇ���I�����m=����n|�#*���C�x���"�ȆU�����
O�v%����4�����M����f��t`*v,"B�Z��NF�̮Q+���i
��fH��rǫo�p1E�[���k�$ΫoY���Q��o���Dh94kR�s�~���K ��G��x�t����J�(}G	�?v
r�^�d�/�lа��`+�$��Q�U��xm�y	$,�H| �yz;@;p����^xI��a�_��^s�_�D�{X��^�1+�[��0PO�>�ep0�;�S�I�e�o���^vj\�RŬno��_p+=��aT�7i���ҩPt8�9h���`�FW�R��,0�9���wn �é�����-Ŏ��P�1�v�[����C��)^����:z�'�_�dH�V��l����^�K*��S�z`�ṙ��8�PQ��	�A`��3{<�(����������v���l��>U�����>L>�sG�.�{�4�V�z��V�;M�
|�§͸��r��K�/��o���M�ד�U��N�����po�_�����4���.���?mR�-^�fױ(����Bk��u>��D,���?�
bY]��F,z�Q⢎��B��D�F���q1�ΣM��+�\h���B����"�ܣ��X�q���oL�.Iܨŗ��ŻS|�7�!�(�g� ��)�I5�ڦ�O��H�X���Zq�u�qA�Q���0Z�
& ��q_j�J뗇�~�AI�a����IY'�"�5a����n�Ϥ������b��~��tCwȞ2�:��S��S��_i�i���@�Jߍ���Y!h��N�7������Y��
���$u+���@�w~W���AT��6S/c���l�"X�Y������R�^�������q�}��&����Uw!:~3���R��B�O*m�'�_�I�Y�Ib�_�T��F����X��@:���O�L�� T~�s�Sw�q1��b��YT��"ԃ��r*�s�)��n�5Cq+V�,����N@I?F<9�lҹ�����t����aJe�D]������|2Uo)sYO�A ��������� F�y�I�I��^"��Ľf���m1 ���q��S�%EUOZGZ��F�;�jkpωP�%`I�M<�	hjy����#ǉş�@m�}���쨊��/��>{�.�/&�7�Ԛ;o�$��� ��,E�T��k~� O`x��J}�f%�����;z�Ol(�j�t�2�|I�} �d4)4մ4�;Q�
I�3��9}'n:aXex]g�d�mNT�qx�����;/eV*�Y��� S���+�C:<�V���.@��Й����������8���W1a���q����_}~��`��>|�6��׎U���FGY�1O��h�VwT݇��ȅ^�b��o�d#Z���0�휳E+�� q� i�C��}���p7/<��]{�+3�F�ȼrG���s'������&��jAH{�߶�G�\2����0�3R|(�b��TsJ��5�Es�c��ir���r�:/�m�y�J�mS�jJ�|c���F�ޚ�xV���;)vE�f�8J�*o_��پ�s�1�)�[͍�DK8��<�*�H<y���W�c����<+�	��a��� 3J��S�(v;��)��I�rL�&�����U�)DT;�%C�%�7��j�����%��9����r�P�e��b+�j�����}x~�șH�&�AK�MP�u�N3tk��R3Y�Y��~��=3.��?c�$Un����������~c�A�qw����F�h*���.]�������z�;���|�P�P������I>]1ӣ���t]J�$K����ᓑ�%*��f�-k�f��H�0-�':Wlf��]+!��u4����ڻ>5�ae�����F�<�͜L��1�o�,��.;��S�~��3�<僦����@����Ly��w*�����Q)2"d�y>��4apG4:
��O���F�� )q�0�̄a,�,��ͦ<�?�A󉟑Dp������oĸ�gLA�>Ȥ�Fl�X���{{J���^��afe��]�	j��l��E��>E����h�ڠ"S��u!���s�*��*��LZ4S��O���݃F�pp�:R��B�E�{�*L|�lQ�}:S��0�{ǂ1����$ XF���ђ$��`�e,ś�Q-�b�bn���S�cFDʼ��ĐE�	��x��wX7`|�����~������Y���Y���i?'����K*O�澕~8᢮��h_�I�h��8>y����e�a��q�.���%ts䅚�VִTb.����v�e�(PbL���^+���[��s4j~N���)����Uś�����x�F�������o'�������[��|%��N4c!������p�0.��ɳT5� �Tb���Ý�'^�A	!Oq����S���鏓V�
܀s���V��D8�P��-�}�����\Չ|�O	P7�g^�_}�a����,��w�E���i��"ˋ����/*�����$���L鄅���#��nm��b�yIb���L��E�������Spmƻ.����5�$��Rb��iA��c������
�Qtw��ʇ���RP��@q�	K_����K�յ�b��H�S솖�̀���N�=:�0D?�.���(V廜����ʁ�a'�j=�1\�j�$�@�l�Q�ݙغ9�lh���l�U�V-�����9���w����/�3���ܰ�!�O	i��a�HE��_��u�#�-E=�����D+���e|�Fw���R�,� C)͡|�X�ǹ��V�zʂ�`����D�퓦:�+hӬ1�����?��E��K͌�W��R�@1�R� �{k��ܼ� �KS-�����Ȥĉ��uZ��1�1�E�
$-�]����ϥ��V�	��1�V��{�JU\��ˑSM��9?�lsw:���6�Z�%�W���	���q�Po=L��ݼw������\']Wq��/��@�%��\�3F�l���$��pHQD���m#��Z;L�n���}/o�}؋�8�ˡ!I��l0�DSuv�\Ϯ�Q(��/���*:��]?B��|���	x|�ꉋ�)���-�|噍�f	�����T�E=�Y���;���3|�v����õ:�R�]7)��y�k�F���1�@K3{%��'2+�0�����~鏏�=�,�&�qkm�Xy���*�r��w$Y�3�������J��]�zFX��?i����a8�X7}yg��ϐ�%L[Yͧ��ˠ@L(1�]R8�}����P8֋��<�7K�����B=	���{��!�ԾD	�ɼǖ����LB2J2���ƻ��:�'�6�;�@-�ncw��♩D� Ӑsʪ��R�:�bCT�Rӛl^��X?��O�U�7�+�x��Y�Î����=S���:�'L���� e��=D�T����s�XT�c2]�]������@V۲͸`�o�U�&�eOy_�D��J"�	4�YaB/�ހ����0el���x�#@���԰�ЃfZv�LS�}�p�	���@ؗ���"t��� �;3Pu{�F#���;��1>���X��@P>N�"��ў�8��&�3�Ej�^�q/��v�پ�gED3�3c%��� p���7Z���o:��	M�m�单��p6ٗ�m������Ð\F�F�-U<e�	�L�{������1����M��;�II� s@����W�g�f��@����'6����qǹ-^}������(q�	�j�P}���̥M�� a�����[ݰ�6�i�ڢ�ƍ~��|�H�޻?�m����.x�Cѵ!og��;]�,
�]���My��Pd���#��Xz��/F��
/�֕��B����^�bcK���&����M�5�4ԩ�*T	��ʼ5no�R^��Z�.��|R��%<^�`>��]U�����P�8�e0J�٦s%��{�t�\��f��J��8��d$*Yu�8��I�%�����6���=X�o
��{�
H���*���)~"&������+z��61�&S(��N�k�b2�k�����
=�*����\̓�v��>�X�y��WrK�f����{��Qq� >��{m�⸆�(�_��ɪ��M�$�aDi£��7<�IZ/��;��\������IAc���L����0ӹ}H�]������|~�Q�M���n�s�y5��N�U�HV��yW�Y�#ݼ��FZ�Q�a�bGd�un���,���I;�X�����0C�&��O���<-E��V�$��
�j�"D�Z�X{,i3��7MS2����C'L����"��Jj�q��8���)*���e�BQ���+s`�/�X2��S*�s����d5nO�-j�Ck��f��$�lE�I��� ��b���S�zE1 _�:�V�����n��#�S6�"
��5)仴Hu�5�~�9���������X��9�+}!vXr,�n�!��N��!��en�����S�l��~��\W+b�?_q��+ܮB9z�X�k���W��I6�v����{��g��Չ���r6�wv���@aũ���8�>G��Ƴ�
��sGs�ѓɜ2�/��G_��E-�?]��4Q;©x	����1�7��80|�%ůg��tbk�?rp�\x={�3+.�Hf�b�4��Qv/{]&�MK�	��r cq(I�9�>��x�J�`!�+u�"�"&����
/�mKkZL42"e��e�,ģB����מ�v����Pߗr���+�~�е��I�w[g�����T3���L�	��<�o�����}gͳc&��R��Ϸw��Z-\���{	���Y�u26q\�^7bBg��E�O�V�)������p�΃����k{j��|�N*N/�+�%��ϓfח;��{m���D5p-�EB�L�j��.{��[�4�M�l܁meĀ}��"b����s�N_�/�_m����a*S�2K�q�/�����R��=�9$�l>9�P]K |-�+S��U4.�1�g�,��-df�]>&�%�{>�W��&Q}@1Y�"�p�S��S��/50P�q�j)�ٍq�w��p��ǚ�#��%�s½��.gҫ-�u�T2ř�窩�,h��ؗ�v�����d��+��}-B	��_-����d䌉��l����\�2�GD��_���Zo7LF�*U+��%3����@�Q~I�(�֤2,����[�����=�U�+k�֗��!Ƅ��"W���"��w�a���5����ӫ�>�b�x���E���>���@J�%���U��	S$��s����:^P']#�<e+�H(��3��Si��DE�Gdo%�����2"i�U3+���.b*��K�bˈ��x[�$�!��U�a�9�����O�V�A����@Zr�Y_���zY}�� pp*Qqm�5WdEO��j�H,�{���+�����u��&Vr��v��倭6j
����$=�,��P�s�7 <�Ѱ[ھStc������Ƀ2"J��9b9d�� 
��%�х�
S���۞Vآk�r�r�������0bt|ȗ?rZi#�_����!�7rW�LZ��ap0���#��=�h���qS&8�r���ۈ^��gOr�	=�g� ��٘�,mƚ�Ke����0g��b���V�4B'xl�-:�Ob%f>�C�+]ƅ��R�ˀ���~��i����v����.13��s��i
�����u�{�Օ��_F;F��4�5Ƚ�&YV�ѻ̕oґ��ں�ѯl�+���'�]�o8��`����f�M��$�٪q�o���C_k��-�o���u�W��R��\*߻�%��!����網�*�!w�]W�	��|(Q$�k��Ŋ��w���e��ŕ�	2đrAz�$.!8>�yN��q��>���]L�:�u^�������:Ԧj\A&�9ьɠu�
�-׮U�{�UG�*ꃶ�D�ĩ��Bެ9��<�2q7�qm�V~���m"�΅q竔	#���H�[z���'�?�
�~�����Vp���8��+�N����T� _v�4J7��qJ�"m�#�B�u�)Ĩ����]�>�^tL>H]I�m�Z�C��ί3��|H�@� ������LZiy4x�l���h�/`UV���.��>�%�ƗY��2�oܬN�o�(\������p���8׽.'�b85S7		�0�L(Fq;&�Ti���C�X��Lj�\�G|��
@�������$��&��������!W��W�q���CD������!���S؄�� �!oM�0��_�qBԑ*�0��+��q��7w���+I0Y���.#��|�KW>O(4���*��l��$`F
?~YP����X���4�t|�@Y&��h���3g��������[d]�ۄ��-�wsZ!�9����<�鬚�,�$�ۭ���8�O��l4ix%f�E�ۢ\0��p�p���
�H�ĺ��n6��D�W7E!�PBJ�����{Teg���K*_=��?t���5�<g_�L&r=m���=���r�On����͗S) iPW%3�#!���/� �z8�}��T�Hu
-��4<��?���o�$�O��U�2j:�)�Y���f�>��*p�)y�HPݮ���oF�|�n���es`�8�ʡw��sWy��a�؎�� �q�ƹ�`��
5D+F�Y6r�N7ui������ʛrxCx����u6u�`�Ii��z7�F?&s�7��Ӹ�n��`@;C��D+'/���K�'z�+5�����@�R�S!2+���v� "egD�ՀC�{No��^�y�	�Idf�hU^��z��S�H�8,1M�%ͯVbO^i�%C�O���2���|]Zo�r�ϱ��R^����M��3%�7p���JƎ�:P����mO����v`P���	���9F/=%�_n��~�䪡͊�1/-V�I����Z����gw��	���˔��P�s[y�S2zç�*�����X�j��9��ӌ�jI��(g^f��>�/�|1ė�{�����7����O����T�d=�=�w��ã+�]$lZ���2����2��g_�BȉE3���{wt!D����d��������.l�!^�s��u�9�b4z�kmZv� �w�- ��6>��;<�`�VDX�|ΌX��|AoJ}V��T�X��ۧ����)��C4��!�;�C���h��j=�44<LU$>�8�O�ܛkBC�|oy,�s_�G״������K��!��]�8,��	 ������]ߒ�y��W5S;Us�̱���9ݽL*F8u
R�c�.H.�h���Y`��=2"���W�,hh�������Z ��BM�-�q���ԡ��<�������ۋ�ݬ`R�o�`���7X�4ނ*�S�`��R;cQ�mB���H��h�{-y�y� 3����jB�]07�)60����%m/BхСTc�ԛ��6�:$�g�|[�Bn�R耠H���:��88�?��i�!�c�ޞ�B�?Z��Ю�A��6X�nˡ,��6�_����&q��󰊂���!��}yC�=F��.-i�#˩��|4G�����0��yRi�?t&妇��:x%O��q&t�i���u�I��i��*T�4��z.7K.�	����Va"�lj�Aɢ0���� bH�Z��h��f5~of~��8�@C���!�N�J�n��Ӻ�w�.~�v��5/���.:�Ա1�Z�+ڠ�?`S�� �v�Cݗ��E:��,�mt-m�R�y"K*���������l�'42����![���T��*�.&�Z����J����������w��b�?���m/m��q��@Y��+��n���'��e'��<��nW�K�Xc�CK��S��}B���.[>�q��gFk�W��#�!#1�ٚC��q�>�;ҽ�Y�ج�E�����2k.>=H��2
vb��*�>7�%��2�	��2@o��fG��7�//%�yGW
r�jW���~T��Jnxoxd0�A�(_�,���ݧ�j����z�ؾEA������h�][��w4 ��}�,��mM���no����ͺ�� ���ď���c�cK�L�w;�ʆ�A�՟���vSʄ8�Z��s��w�]��>.>;b��U��v��n`��-�zac/QJ�|�1��E>Ԗeu��%���=�."Jun=,U���[B��U繺�έ}\��_�l��n�d�u�(�8�5aپ^�ͤ�W8�e�Ü5�G����$'R��Ow��u>��ñ�z��ng��k�g��<�T���}HWpu�wJ$���:q��tBe�]v�9W� У�}-l���Gcُ ��H�������[���9�X亝�����u��V�Zy�
��	P�^�l��RB:�BuF�� ᕆ�H����~����ʞ��p�-Q��M��'H�)���d.�s~���?�R`���>���Q�@o��x�`E}P�.�iu�ab�+&3������݄z㢪��qX�F��!��Q��;��4�O��Tߙ�M���=r�O��)l���~� �.s/�?��ݓ��G���r��x�7��`�شc�_�M�i%�d˄i��:\2s�� $��sڎη����B�����<��I�����W�/����v��6����.1�:'N�1�Vڷ!�o�b��͆5���� a<E��S0[�&x~P5V��Q��غ�zO�zN�TE�qcVݯca���f�Zb�(�)�a��&�]���V1lVg)�W����V����aVcT�5U�ֺ��6�E�F�F���2E�HJ��IWx
3aT���ڞ�fvQS����3/����u<kH�x,��e׮�x�T$��Fu�j��Q�lȘoW��R�%�s��`�VyH�>%M���I�WD`ty��]E k*G��%q׼e��T���Shw����av�8�>h۽R=��^��H�~�2�B�b��a˽�?ˍ?k����@�O��\�m"�p�oz����=)4(L}���[�5�gmm�h�Ehr���l��> �M�s�����h���d��!����I�P���f�B4)g_s�����H7!��E]�b�O8<?3xM��]_<3���	#����h�,Nk6]5'0�MzU�����/'����},�˧��O�D1Vw��͵�G��8��)#�Ѳ; �5�� ���^�'����"��%�o~&��լ��yyEmA#e*�1��h����|�B�{`eM�J*Y/F���tis~*_
�J�~�l&���=��Q̂��
�[����Q�u�(cL�{'���$�wġ���n�.� �2�pZ	��Y�P�r����N����-�*�\��d�/q��om(��F��J��/�Nz�=�-YtT4��?L�`&Ҙ1Z�o�N�n��:dr�������2�)���5�&f�N�2�� �*e`c)���AY'����A��Nt�R-�_{	i����X6_��G����,`�3�[�c?��SF�}�Sà@���&���PF"g����޳�ͺc# V�ި.�?m���8�ڦFed8>'H�]�]^��D%ㄏ.��բ�rK�|�`�g��e��9r��ӑ��2��C.��XS���Bb)�f&����8L$4�$B��O��S������s$6��N+%k
m�+/����:Ӱ�*- Ã�x�q�pZ�4q*��;�M���ۭlTCL��D'�r�7�9<3�}O�C���ዖ�9O��:]�k	�Vj���m��� &'��wsW�"���Z��R�.����]����ިU7_S��l5��7Z�'ⓛ�!���}���C��?�Iz��?v �#l���beܐ��p���)hoO!�l��7л��E2c��w��=عe�
���=�C�`�s��dl��=�ҷ0Pt�^b��>�"f|u�69�Ÿ}�(l���?��K������HN��;��[�׊�Q����yB}���ˍ/�;t+��4��|L6o%���,���S\��v�!��I���Ēb.ø!��*�O�ڹ�E5���-.[ٌ��ܼ���蜮?�]�>�5�(��EY��X�l%���x|6�X�c���|���T&�0M}@����7��6�R.���6u$UZ��d�7Ok!�w��2��5��E�##m�Z� ���FkK y�]O7���E�Ո�@�B��:�]tR�@]�6�"҃C���$����`-��yj�ɿm����~ݛ��������hi�a�2�T_�^��Y�������䯂t�顷AA5I[�mb����� ����� �	~��'z�X-̺�n���N-)ٚ/�A�s�������?��q6tp����($t�ǲ��&���eN!P�6�M���xO@�8�$qd�����`h�o
LڜϮD��3+�b�����w;�f���3���ċdݢ��R?��K>�&nG���b�*l��Yi���Zj�龾p8�����7��I|�����*��J)/�B�F_��{��2M��v}�H�@�
�iir�<��h�<��AT�K�x�-g:z���Rtx"�5��
~>�vnco_�5&����xDs/��$h���F\�΅y������5!�6X6�>5�(
�/����u��҉	E���~�rB>"!���E9����G+L�f�KDII�Ҝ�g��q�o0��*?u=翆�H��[��V?�I��s��u���?Rq��&�J)��H���T�-�8.eo]t7���9|sbb�L)�����'�N|�e�M����؎����K��D�a��<m�L|�)瘈!�+_U=�@�QѴ�"P��q�;u-{�_�u���m��h�[��eR������U��a��L�u�p�/3I��3le��RFZ��rR�4q7�c?���w�8T�˵L�~�@�������5l>�&]��|U�-k�ou�On]%Dm�c#�^�u�>�4��i�p�����Z�#�]���$_`h�J�ց�_�q|a���������p�<�<H��eC]��xdW.�3G9�èŌK��8eO��>i%�+��q��Ѳ*��8��9��%���`���{Qݙ��f\�T����1^���>m��h=�J����b�y ��s3�į���>���αw�q�d�)��-|�A�d�e=s���SZb������Mt_�H� 1j�{�����յ�Н�Я`qMD�}+����d�d�^1�@����������|�q�u����V�S䨼�;��&�,��?~4Q��_g�q@y&zb�L�Y�<���g���#GuE��������i�	�*S�����٨)(�wz��'nB'w]�n��$��5��	�0��‍0��O�����1s�?-P�>�.E��E�XqNL�=�'/㍵�qW�qt���Q����a�������$�3�4�ټu)����b%l�K�+V޾�&�g�6n]ַ�ӳ�1��U�����qE���?���������@��(����u����2�'cvZ9�/�R7���*�f���"JI�����#>];�/�>�o���^q�)D�J����mO��/K?�^�i��4"���d����u�Ҡ���--�NE����[Y�,��{a5��V?�p��]�eV�������M=�o�L0����+~�O�z�5Y���\��"�������ֶ���3_�g��qi<���gC�v�s�$�qM���3�T���R)��J&��w	�G�`�7����R<��N��ݤ#;ɪ�&��j<lB���Ƚ�	H��y��|"�t�qh8NHA}#ϙ�Z/Q5�{6Y��Aިǫ7Y�l�H��:��d����K
I� s}+w�4#���"��c�*>>�G��}n��`���"��A��B:���PO�H��)��M0� cQm��X�v���5�N���Ȝ��H!k�2�vr�A��ϊ�?�\~�ow���W�pD:�}��p���u=ꍇ�h���TAA�$��P}oR�յ���^�,�����
`��������s�Ը����ټ��!M�}q�����[xAG�Z���s �V�/�˗�?{�}s�'fOSTm�%���jeJ���
p����	N,�����ʛSaХӉ�@D���(���SE�{�R�˹��7cb;�`.�_��Eڕ��B�����ҽV�{���Zw-��;��Ƶ�F�v�ݟ&|��֕��(T�J(�&,B�d2�H���eJ���6PR��1���^���H��Mt9R馀�G�WqұS����yr�Y�@�x�c�G�<�+� �P\T���7G����B��<qC��}�~ۍ-$����_;�\��Y��>�J!�B��h�ge��Tj��o����+ϒ���K���sOA�M��b�߇� �i��x�
�	����X��
3NA��XC�"�ˊl�z��W>�@����J�R�`��㟁��z��T<ҷ@��v�bM#�s�	^q�FA�ߘ?x����6���ո�͢�1<�d���|���'z�ۤ++�����~������� (�+�r�~�T:�X�tc�R��ݫ`M�]�ao�-ɵ�)�&jO�W`�֞�!0��v�(��kWCJ���M�����W��f�Y�uw�R�5��нs�^�Q�{�X^-y��1c$�?�ר�E�a!$0��q�Y���A=.�����G2*��5���ټr�D{|=h��v"�&��_g{��׏x��jF`��>c��8�ς�d�{���_oC���u�U���s�`!^Ǣ�b�������r�P�컑�߶�&cG綥hyT�m`\+�_����kj����Gb�䭭=RAj�h�?u���	������s�:Y��\J9�n�L��q2����Ao����_��}�����Z�)�iU���` a�����_�S��k�^ƪ�Jf>��6yN=��5l�@{w���Bli���3�q$Ė�	壡��k��x�����e~�~�Wji.r��`��f5V��O�� OO��Fw�~�P��'6T�5`C���x������~�*0va�౛bjL`) rXJ�T�ᬬ�=X��0Y��R��b��B�c�h8�35���w~H���<"���2,�����LQs��W/s����� Q��¼�"�y	Jh'�:�}F@���)�}ʫ���Z���-X5�vm	+��"k��eVO��w`�'M���栁����|�X{�o�t�0g*ѵ�����/ �M�V��@�T3ʱ"W�N/d`N}��)S�K�{��E����e
����Xg,P'e�#���u��K�$�,뫤�?�����D�Z���|�|D+�,K׻F�%�Q�.+C�8��	�#�+8݈�v�P2x��~t��"�đ,릣:E2���)H�1�"`#Ĺ�U�u!��}��=�,;B��H���?͘�Ș�x�D@޹��k��G�c�۸V_��d��`p>��sX�����eLK/�kˑ1;�Lۯn��:g^-�����ﱦ8��F�4���\ �����?w�D6�w_\�1�pk��K~��'��t_��\&X�n�:	�x�b5�b�~�Fx�V6a҉���������d�� ?�FvU��x+d���H�f���&�_g��/v
���TkX��[F�z��!iu�}�*f"���6��{~���ȓQƧ4���a|!�o�E]2U�+.����+W�|��/�٥�yi�1�>��ނ�$�?�ῄY�G� �Gb�����6G%\�ޔ�k�OX�[�m}��p{�+I�����"�^'$;xl��%a�h�#0�X�I|�/��]�G��A١��(Q���-eEBm8�-��|o����2@��|�.�ɠ������T,h�18#��\�9Az�x�N�4�Ě�[�;2����}b<x� /��^���i�M�>��2�ȶ����6�)�e���ɯΝ=N��%��{���Z���NT�d��6������@�z�E'Wo�ъ�A��3�y�a��	�E�Of�Ѐ��� �����Ȅ�ٸ�P��^Gb�$��Yj�W�ҷ؅j����k��U��د�g��3C��G�A(�~9�^��Z�6����I���o�)>[��3�gr4c�@��je[�;�©���?�ى���p��IR3z�-{���R}�ۻ��م���vfMg�z��ގyP�os޺��o����?i�F��|v� �E�@w=y���zR1�S��t�J�6�0=%]`�N�;a�0J�c�+�����=)�?őw�I�>���0����$���Y����r�-�i(��{^mla��я��o^n>����&�U�`��h��ݶl��*݇lj%�(f�����#B�ѡ�d 澿}���S���6k�r��=�v�L�	 <+�M���J�m�:��FO�u-�II�߿��voc��MY�O����cIN1�t��0���I�\@gό;��O����c
�����1�D�J�Z�
�H1���_[��W8w\)&|ϳV������}<���.LP����=�Czc�`L]ب���%U��r���~Z� ��qC�]	Ɏ�>8⻞�[�"���-���F��x���	B'���e�am>1r:���k#���?�'�q��o(��q��w��^O��$��~Π�Y�72�d� ��`�=��U��γ!�N�E�N�F9�����"p�޼�(�C������e�؂Di�l>�xi�A� �.w~�z�`bG��OD���r��{�`x]��{�4Q@�sJ���΂���Xq,T���1�FĬf�o$�Ԩ�>FI�o�n���Ƈ�.�τ]�����ƌ&��]�E�iu�c)�ij�N�oJ.*$�EK��ju��e|�ؒ{��'��~��������co�p7�A�XA���������Ĵ��s�G+�/mth��g�w
>���I��>��)��J��wbqb9�")1�K�R����2>`��H �l&�h�u�(��R�B�P�4��@/�Z���AS1۝�?LPU���*4�b��wQ��y{C.�oc�-��dH<[�rP��hF���F?��	X�9*��>�RP:f�e�z�T�Mn�����#ҥ������T��f��}���oAt��qף�@bb_��$Օ�	Ĳz�u�&`ėח��7�D6��!�����W���oo����_=�ll]�F��m��ӆx8��^�����v�UQ�� ���I�_���	��U,���K)¿��m��2��5��y��@ܽZ��F�:"��s
%n�NQ]���\��2�X� X����ý��n�K��f4щƿ�f��U�����Ņ�iLN3��i����ڏl�r���	�h�[x^cH��JL��^�h�����t�d2�nJ!��TwK*t�7�����9Z!�P(�Zǲ˦A���3�W��s�i
w��5�N�ǟg�� c�Q5ǂj���KmgΓ�_~��9�����#m�[�%� ���G`b�u�����/XҜsޮ��b��+�xB&��B��J��C�2kٲG/G�&���q�4�`q^\d80�wA� 7�0Wۉm��N�g��oA&v��?[a=~:���Y���L?hY�T�V�'Ö�T��W�"�۲J�@J�IRd-��u�Z������$�PIT(����HV,A �ܩ�Q)�2�!�J#��Tڟ`��Quxh �(��LO�s)݋�?�OA>��۴�K��0��b�T�Ϲ"hM�(�q����O��pXC��A@�3�y�/���_�{���S��I�ZA�O
����"@z@��SS;��&G���'�U��*z"y�_V�X��ڌ+��T���k%9ϓ)8(4��S	��5&�� �N2��?��?0�8K��g}��,��HM�M���P<�쮵�zG����vG������64�!�.ۓyr�r���Z�W�P��?����7�Q`�/p����%��S��+���+�?��$��#|�򯰜$��������t��V�i�е�$_=X�^���S�D�L��H׎K��Տ����;b;���^� ��>�_��~z���!2�̝���G/�y��:|� �Gw[��<�M��h�4��Y����,c_���YȮ+�ꌢ����L�l 믬'�����Nr
�֍��k4?/���P�dhw?uj}Y��M��"�_�r?Ee.N��L�=?T�^��v�r#��8��=�=~$�a��S61�et�$O��_r���y]�ڀy��o����ﰩS�/|��Ĩ��Z]v���}-=�a�t
�5ձ���ԵxY�vl��.�_�����[4�V0f��v�8��֟����/'#�~L���Tf�G�{�ec�!P8�Q�����Y���B��O��,pE�����"�N壊6��65�$6{�~�2�l���c>�4^��(¢�_��+����ާ!\�d(�u�Yʃ��Ť�r%&P���� �zȰ?��َ\�uϴ﷝�� EsJlQ˷���/o��5'����P��6=��2ZrT��>�8Y��x� Ɠ_��e&�'�/2����,d����̝d`5����a��n)�ї��-��،g��P���k.+(P���?5qn�~�dc�N�].Gc�c����T�L�������%�\��
�T6m����arC9��\:P��.z{��s�tp �����	
u�ϵ����d8�� ?�K��b����9�w�]
�
�8��'7�a��C(L��8��,�u����f �T�9m�]?;d�F�&�4'��cf�_$)N��-��d���l#jat~�j.�JןM\�~�����/��1�� ��b3�8�T$a|)s��:쇅�DD�Xb���?���L4sAh�*?�����>Pm&\�����ϐf:VM�G��22T��rը@�M A*պҝԕ�6;�'��+��T Z2���-Ѓ_�Z���������K�M+�Q����C!Z�؝���Č�Y?�����h�Uk:����S�`T��G��yl�4^�X�?޻v��7�F���i�����${�K�,�m��,�#t�����s% ���W���C�O���HJ��B���q�����$�~�,g�,a8���-P'��F���Fd�W"��4+�r��/��%���� ����BWh
w#�BJ ���􂣭�͟��:��.�X�#��>-���?�=w���)\�͒x~tڂ1�'&�䖠2��U]bհ���c�+�M�q� N`�:WVRϪ��w����8N��2nd`R�E�,Y;�e^�&%F	5{��'S�J(���S~E�-K�c3w��I�g]*`���"�o֧��kO���5:�$#����	�a�"׏"����ͦ�O�� �Y4(�oPi,�W��.A������-S�k���g,)G 1_x��~3���� `���7��a5�����F��,�	�ˤn-�j�TO�
_�S=�G��$��N�F�A{�h�<��<��<q��F����\(o���ܸ�d��&W��uE���?V(T4 �vJ�=�?�=���@�&���|9��5J8*-2#m4���e���9��r�6���C`@g�OG-t'K��l��E����]0� ��4M�c�W���y�J08�2s#<�3|@���8�>�vF[�0׽[uh�NX�p��_�I�d�U@���W8��x���d�#��Y�S�p��-NQkh|)�U�MJ�J�RR��k `��"�^����㲲8B����JB���BL��m�X��o�B�!�ϑz����1�!M������͗%���Xur���-�:��J��|�]�u�T��b8}��}Z�7��߲��Ĵya��T��_�̘8��ӎLÅ�!�S��*�?���}ǳV�Q���~�P��K:W�b���o������j�ځ[Mq��-ݝ��8��S���+�U{g�Qr��v���r�N��zsw�[��yid�\�.�X��S�L;��'˘LQY���{r� ������,�LJ�	x3�0]R%iX ږ��Y]�%λ�8{̍��)�E��*�����Ч���+�K�m
DZ�-D��䬅w���|ӎ��8�b�0.�,�~1Ȥ.%e�A]��e���
��%�Ai7�g$XU��s+��~�( 9Ѹ�嵔;��� �Jm��j��J�MH��*ч��%^s�F	��8
���Gen�܍�l#I-JHy�Ⱦo'�J�'<���h�����rNj,-��{��A�do��L=��bT�?�Y��FO0��������~͐�<a9����6��oTPǚ�%�V�h0	p�� �
�1ʉ��ƶ�x"o`C�|��Zs�'6W���D~�ެo�NfD��X���_�0�w�ظ��V���{U8i
�ٗ��idn��xG�2{_��,��A�:c�Rx"wo5S�E��k&��.]�����f:,WG���4�A����)�꽣и,ݐ� ���G���(u������������F�����I�!E��{3=T�>���X�9K�b-w��Z��b?L�)�׀�KI��>Hkph�7��DSl��u1��nv�z�����$�;E8��f0㚌	၈VB��z�0	0^�RZ�_>B&���5y8M���Àl���&$F �� ��}1�Dx�&�Y�P~��P�L�#Q�������;�}�4��>�;�~���&Mwe�ܐ�ˏ52��U�D�@�;�u�'F_U��Xq샗Bt�3X;�Yݖ`:� 0��~��	��0�q`�V�����BŚ�3�+�F��H*L[_Pu�}?79�~��lo�xL+�q}�L�P7��A���\����sl���T��jv�����V��C��{���|O��*�y|f�V�������\6�z��j�1q�V����K��x�˚� �frQ��.7|�éoP��Nv�^��o:/	Rp'��w���".�DV��J�5r����/,��(ܢ'� �ۍ�ּ�0�Y�߄y��#uR`#g���G�~W����p�e��Â����J�GM/��A�P��^�l%Y@����i3/L��ݼ7�R����z����<R,}]3��K1xF1\I��Be�~�+͔��j@=+�Ϳ:���g��-��c>�t��~]U]�؄��9���/���vt�_��M���i.D͊d����T��7ܖ����<����
W�����s��As2Y ��vOQ=��m�>�)u�����u���+�mw�:0��sR�����n���V.�A��r&P����4�8Ws��o��3s�Q5�n�@X�:J�ac^������~�@� �j��`Y��'���__4ʠ6�[]���z-%wD��1XI����|}�HҬ �,�=\|Ǽ|����J-���,	��B�����_�@U���3�'"�$�,F�`�)7��1Q����$�����������}�"β�E�V�@�u��-Yф��q�mk $5$�1�H2���}Ԥ�I�$x�pq�2Bt/J�^�j\����S Xj�M��g$�G
U4@�S� �>��%�������g����� ���T[�lD�j��Su��~���P���Pq����9=�uIFqj"��mk��T׌;�1��	ٞ:�f��Z ;����B�a/V#���yZИ�=��\3���3�5�J�)H��^Y)��wLg~�T���(>||G�hʼ!l�H�d��1<����G�����~���X\1h��	�FV��CiF���dD�ђ�D7��(�H�����X����E��CY�ċ�QMi�0��:���	C�|.��ap��vj��t~���Ph�l"�.k�E|��4�k����_�`�� մ�wd�Eg�#r�e���d��<��dֵ�����ǲ@�jP������x���^�QF4��*��k"��~Mh֏j,˴e����
�-��?u.c .r$�Y���_IL3l2��r?����-��
�u`c8¤,� trW�\6�²�]R�\hf4;�"�.�1�����*����s���ІM���\�@��{N?��	�n�~����������������}(M��rj�h���[US[U�H��I�b�(h�mM�WN�	��ɜPC��94}g"}�Q��#v�ߟ�
�����8ߍh�}E1@��(��J�'
W��t(����v��R��<^ûG*���2�n��{�6�g&Nr���A
�D<��?��^xBp#� �Ҝ�a`�����2DTl������������j5��xq�ؼ�̷-�|d#�'�W���pw7�Q��j]8��y�HxR����o��վ�,���QUSN�0l3Q��']�ٴ�S��O����^5�W���t:7�fĨw<i��<4I�d��S�������"�bp)X�S
9a-m�C:�l��r@|�F��㫑�c���i:ib~r���n����3Y��&�Cʓ�-��7P�x�2o��31�U����\-��m`���'���	�:��#u�
��q	ń����$T�ЇN�~7b+���������V�f��CD����(��Nk;�U�KQº �����4�9�&�M��M#���_�i�����Y��qƳ�`*�w~ ��`�aBU
��=Mqk�A��`E���oM�J��GKO�fFj�&wb+Պ	Y
T&�Ƈ�=�D��[)�	7ad/��R�7�����i�m3����쳽P��R#���tC�@v��w�	�^�TX�V�H6�OV>G���͋�@7�5�U��EZOխ{��Y�Hek���0:{�p��&�_^ �鐸���>��$&KjG|X-��@�>h�[�����M x\0S���1X���vV��� �V'�����6�![�h$ ������V��r�/���~`�G�p{{^2��Y�:!Kr}��	��5�7J�e1�q��>����`��|좡8��jp�QQ^^���#��?� �����_��;�ԙ?��.T�2����B�$����\�}������q��FT<w�ɎU>f���%�f�)m�i9��vk3��eti�FE0šLbY��o��*#,�t�`K�����w�E�(�0>����9}W\����� ��P�"C��c\f�'Q�v�������BBWC:�6�>�{��͠�Þ�Wj1�G�q�鮓ݯC+�im� �Q �ZD��:���u~��عA_��$���myg]`l꧑`	F��VAz�����5���M1��9r�F�貃��.Ã9YB�IT
�]�:�?Yk��):=x�[�$k�@�-������0�z�e$U��mz�uFOZ.����L��цH�c�ľ�!����DxB�2��[1��`��>'�[�h�Ǚ�ȗ`���3�~��Z��W��6������̘��H�H����:�8-M�j/H���]��;n3�!�q?�>�Z͋���������MP/P�p�񬿧J8���G��X�q�����@�Ӌ���g{�Ȁ�.4}�X�5'#�{'�c�F����t=Ʈ�Vŕ��9�<h�?���IZ4S�ƀ�]�g��m9�&���9d|��R�+�Q�������WG1�41s�[o���j�*z��WD��
Ǹ!�	�<�������Г10@��Ƣ ��8��Zl���X�O#�V2����ψ�)f�h�2X����q,��ѱ���B����hWR�i�9��]������3��ױ$9(Չ)Zl�E���p���p���0a��&��S��o��!&���H��#=�6d�ypc-;F�W����I�I|+E�K��I�m-J|0|rW8��7'*S�>i�J9?��/o��B5�U�z����1��+tq��|M�T}{��b�"�*|^8�:���c�����O�JE�U܀�0�t}.�K�#�,��Ä��v�z���e�-^'z[��b+���N3�X��l�>;�EKK�GV�'�|Vq����(��َW��:�P��v$��,ҫ��mz�|�:U�4ZY6d��̫�d��G���2F&x폧����"��{������=l���vVoWO�Di�ÿU.�g�/�Jaȴ9s�4�!� ��y���A�zYy�0RRl��X�p9�|_h�J��E�&�ǧ��eRu��EK�TT�t<�=��(:j�Dq'N�#`�< ����4�n�j�R��E'Y��^�
:�y��{�����$&'p�+��O��X:���H�a�\3�;x�w�,|1��\��Hr��qA��������v��*��e�$j4ï���}���b�>����^n�"�����F�<t=����шQ��������.���=]���`��=�PP��W��(Ğ�]r���en��Q l���̵�����3G����w��Rq9�K�����}�UAxg?���a?�U!��k��<�A�S�?*� /-�:k�G�� 8&"&K���۾�˞;���"�/;��m�!��?tT2��y���*��`I��߅6@C�v��X�ڭ]�Ş�|�,��L�Ҿ����m]'ŝ�B�ͧ)����5~�|��{�1�{��!���u��ʽ�jr�U[�����l�,rE�v���r��gѨ���	�vkcW���~T�fz�hN-�m�7�Q)*0q�w'�`Q(���\3@�J�-[�僽lNM��4b�ߍ�#W��vf �1��q����G��uO\V ��5u�����6v�ǰ�W��l���W�t@��24m���-cS+qh��kܾ��ŋ�����	L�^�~B�.�b �5)�帑�>�>,���MK��C��|#��,V�A@%~Q/�3�׃A�\A-Y�?Z��R�,f�{��@��0>Y*�w�CŅ���1�T���U��������F0Ta��q��ʍ�o�����	�9R<���6��?��܄Gh4���0p+��������o?Y�A�T!�\�S�z�;ÕW*<�1l�����������Y��GS���~�<o�Q�0�R�f`/I~#����_�A�9�S=ROޯ��}s'ǱZ�ة��9Q�=�]i����O�E~��QK�i�W�-]��D�9Q���Ev��K .C�J����Z5�
C�%��x�(�����@����+g������ֿ�C�bB�z�+�a͟��18Ioa�a�{b�OJ��/_��)�p��x���q_���)�D���H�*�Fģ(��n��:��=H���u� �;�T����Mk�^&n��������	]���ع)�e���[�_;G��1W� +5�Q3}ڗ�r����XK��c�?DT���i���7nUoi�I�R�2���q�%	J�J�|��Tߐ�C�it�>V��dB�8�έ��y������S�L �.o2&^�(OG�v�(��eM��~�87ݿ�������5�i��2��n�g͑ ���;�ҁP��e��R��x����`�P�0�6Lt�-�Lt$�M���*,���ݦ�.�f9��\cƥ�{}]�ߜ�w:�u���Uڙ�R�8YY��M��v&:n�]���M�&��4��?p�Q��D�?��x�>�#}}Xo�mAN�1�#X��/j2�F�,�ʃO\��t��TJUe�u	���q���Pj��UOG�%�&�#?�*�]J�cWM/;e��.@�Á�gM����Y�N`95��	Wy�ܔ�:��	Y��&u�1y߃{J�'�2�O;4c��U�Ų�)p��B��驅���#��-�E��L3�M�{nñxQzz��˕��_����[`R`�� &U=1��S{�R�fc�9b_Ioo3�H�\�־��u�o��8��Jk&�;��L�-{R���<�[%;���?��9<���zc�q6j��6��m�vۘ��ƶm�jؠy7�������d��[�>g��Y��D���&R^��W� �B?R+l�Ð�w�u�a��Uֆ�X��f1���j�T� l�l���	��ʉ��4i��c�E��l+�)@�]V��r�.�.��3������:ibDtm*2ڷW�:�}��Q���lQe��Wy���˽��x�ώ���_4Q�(n�3���:���]�	W�|m_8v����"�I�>�;N�e� �V=��O}�=3X!���F�P�@MO;�@?�l���:�5y�Q%�ڏW���Oi�S�ZO��ɦ��R�ߨB y���j_+8�*�juLrj�5[�zԆ�퉵S0mޤ�Tj�C�vQ�\��������;�FŌlv��W��+%��t��_�������������W4�t8�-�L��P�!� X@�r {�2ב���v������yĘ����o���!]Z��~vD���F,��FN÷�$|��-�>$RZ�~��H�w�4fb��OD6'�Z�Zj?��@`�jk|��������8��f�{zNd�2�������E��{�ȁ_���Zč����~ =��/;uz��1�Ķ�9=V�I9���29Q�)7�J���7��2������ܨ�/��,�'�-��$k5 )4���?[h�=sk�yK��S��B?-��+R��wi��%��;��x���.��\�7,��Z*'ޟ�*o��,�1�2x� �W�4�:Hws_K�$��;����L��	��yK��v�S���չ���I��HZ�(�i��Ռ���W¾�_h/�#x���D��T�}�ǽs����苼~�>j���P�)���A�v��r���y�Jj�&5v<�0[ۍ����p�_����W�-m��9t���5>ˣ�"��X�;B������wE��w}ǽ�mŶv�8�4���f�6h�-��T����Z'�qJ7�,�s%3�S-@�wP��~~]�^�&e}�2<8X�;��	{AP	����/��=����Z�j�f����Oz�M���~s$@�~KA�Eψ�ɯ��`7��7�Y ��N�j����� 3���T����ᖻ�"|�x�DR�
�hr>��tG�DI�8d���	!u���+��Ȱ�8�U½)8A,}�W�Y����;h��5���aP�� ������+pYS���c��
���Mg]?��o<�����-�3���������T�V��k�+e��Ӎ�J���_�������ޔ�@)6�'ً����j��� 	�ɫ ����CN	��+�R$�.��7�{��������}F�׺����7�����u�����C�fZ��3*��Ʒ��*wO�Dw��v��
��� �8���i���J���]�{~ m��y�,���� �`2�O3`c�
�vsO���&�b^�=VmG��'��QǹߢQnS[Z��,��!M	��n;i��C�k��i_m�myG� J%K���w;��K7X��3я"���Z|�_(�x�M����3����uZ�v]�%��@�J�T"����,�!�,+����K���u/-*���t*��a%ޟ�J�[�v*r�G:/]bk��i���O�6zLiM�V�����t�4�mG!���Ԕ������_3-T'==;�Ϡ��%"��R��Ǹ��V�P��!��>�u�FS��bi�������}�k�y����u�z��yv�y�F��+j5tn[�2��Ea�n�,������3<N:Z�O8�\��z��_��KL��9/C8�/OCt�|H���t�)0k�e��r
\��_��?Ԗ؟���*�,�A�nz���y��� £�ص8��{Z\�����-�(���ӿ����d�Z���7����j��f,^`ÇL�u�2g!"����n��� v�^g�)cN�R3�V��C�/G��>!�A��A�z��+��1���ȿ��,a��CEC�^po����3�~��c�+�[�.�������͐H�u�ߘ~��X�#�
��Q�� ꭭����%D廧�r�7mSg����J�����A�t4���˂����^��Q�J����ӓ����;���fBٛ~��I֛��"�E=6X��~������m���;�Nk:�bt�[!{눛�T�R�����`9�h���,B�̻��|ғ]��;�/+���=R�cI�x�o� ����a+f%t@�;U���/�S�WTo�L����(����ٹ���N���[9˯�}������R!�?ɩ7�����-��{/�z\�/K�|��X��}	��eT���{搑�P������E�9u��]w�r7,C�Eqn�PLj���Gh�����x���Q��BxUVZ?�3���_\�ϭ!rT��'!���ż�������rY��у+��7��iyx�T3#�ӗ�o	��󰍜،�H��J�p2�W�/���P�x���ޏ(/M ��O��R���z9�� u�~���u�>������AK-p)n��-����t����6��sj������.:���*<�r�B���@V3�����4<���㺪����ʒ��m�H����O�	��u�� j?�J�|Y����`�l{{,��	<�U�!�&���RWKI�;���<�6����x�ʹ̎�ڂRK~f���;��s�a-d�y|3ל1�S���{�^�z0WΔm|\h�г��p���!��Wpat�P�ӭ�����~�][$������Hf�]�θ�M�-�}�Cw�J��e�;Uk��j�e(�
#�����Fm̧@c����=|�5ՙ�X��n�^���Zs:�W������jk3��ݷNp���~�f�<��5%X����a3�6�-�O������_��������I�f'-�a�r�j��a�B�x(Ե�5�~�'�Na��aG�6L<�M�N�O�{b�`VY���@�郟�V|���/�pѥ(�P6ђ����9������`R	T��/��स#��q�Z�B���9����ONp�^�O؈f����@�j�3{��HE-iL"!S�̫l�bס}�V6��3�ڮ��Sm:�VK�0�a.������<nI���M�Ӓ�f����sz.�����'U�y=�$-�� T:�.|0:qwbMN���Î�4��������y�g/X��������)����S> �@�.*p1�Z��C�%}�\I���Ѽ���;u{|e�U�ǶyÞ&u���)����F�m�IQ`�J1G� ����-�=?pK1���❮
K,)Ӂ�Vף	���������VR>�Z��n���mK�C:�g���}*ըz��9�@��̏Ef0��1_��1�j�.V���{�U�Ǫ{'�~V�nt��]���-� 5��ݒcm:s������~V�}3���f�؍�<y����Dy4�B9T|��Ҽ����69qOu:}�c*������G#P�9dRv�z�W�
jLY�$�6�RRR�?-_<�8���<��Ԍ��M)��o�K��l�N0�GtW��[`ќ�7�<*�"Bt�}�_��=��I;h�����Zlnd�@��	��r+*�د5���V_V7,a�>�^u0 ~Ճ�;^���e�]�q���������gϦW`��^�'�J!�Q��Q��UBV���&еD�r�P�����<'=~����cS�n�E�]h����C����B̊I^�P��[n��x�p\�b_�
��kcz|q���`O���X��e��E���E�iRw�U�}
7�5��Eu�é�n���0d�^�g�{G���-4�;!%̈́؞,2V�J���N&iPv�'�扥 �HD'��J�������){��W<��^��f�L����@�m?�1^�9:�~�����I6�;�\ai3o;//�k�,4�	���_֮��q�5���!66H�)�e��}۹�&N�^ڐ��_�u-���"�� #k����tß����,��醡�l�{O��}-�W�\��%�H���qk��À��Ο:���fB�ą����� �v�=3M軎/]/j�G��95r���t?%��{`�/c��&i����Ssc[,�(�k�%��؄�����MD 	���LL�9����q��]���������m3t�_.�[�j.�,B�X�Ł�����N�s��׼�y�)ׂ���E��Q�V�Թ_�=���&�r�fZb��Q:Z�� s��e;� �Ju���RPz�<��=r�ֆ���s�w?����-8�����Z�M�?e�����RdU��-�~ߣ�gs	(��t!��=g!�V��%SY�G3,=|�6X�>{��dSn�D��WNO��8�|g���qO�j��
UK
K\���V��G�q#�F_ �ߞЫ�4�
���{�*]�(�'�Rz�gqW���w��o��-�̉
�$�op��jp�%l�E*ްx�Er�\�=�J��"�����3��=B�F:�ʠ��粺��b��B'Zo��6�Q��{��.��%�	<mLZ��)w�@�_j~�P��W�l�Ѓ:Zq�+���.X�=�)��\�4O�ŋ�C�w/�4��,�y��j�7�M��.��>�x(y�e���o�	y�֛	GL:bt�s-����eM�Ġ�.�*p
�&g�	�h󳙶�{�ܠU�N�����7o��݇�����jOW�1��J�Kx/�����o�Ÿ"T$���Q`�C�`�̘���-j�%�`z��P�y�$�� t3��]ʜa����}�RT�E��2#C�Z���Z���˪s�ථN�:�(�~�,.s^or��o���_A$�z���+�S�N�����|�6Ƹ�� �]�zx/`�
�~����1iU5=�+����\��vbzS�_��a��f��ʠu%�8��ӏ~L��y[����9��z����I����)_��v�:������}�a��!�b��P�Gk�ބ$��ţ����%����
��f����b��w=NVa�2��Ȼ�9��v�ѵ ��ng%�r*��ղf��2k��/Dܷ̬���F��|&�ِa�B�n�}���\��8ƪ}����m3J�K�,�
T�<���Rv�K�e]&hS�_&Y��ś^r4+�{�B���?zХ���7ƅ�Z�B�P�n�f3/�1��b?>���P;h�2QY^�]�4rϱh��7�)�S3�v��<Bew���sm���S4�|�f�Vv	�^Z�ؽ�}�����5�~�_yݺ��la��)�D?�WD���9��l:��Mp����B�%���yA0ى��~�`��дV��A��a?9�C����8�I��҇섩��O�'ߺ\�|A�h	�g�ig�O'n��\��k��U�-�{O����Ll._ֈ$� �����n`�\c��^�`�_	��;K�Z�%�*4�B��+�FH��'�z9Ga7�T�e�J` �:9[��*�^��%<5�S��(���3k>$1{Rl$<˻�[�m���<�{�E��sdU쎱:�T�&5ڭ��c�s���9��;�p'��	�~O����#V�+���h��@qm��K�����8�̻�3�`B�{��%UG!�F�Ėee����^�~ס����N,�H����͒���/�,eLx�%�[蓼謚f��D�^�ƿ)�G��i�dϙ����E�y@��ʅ;XI�V�wj)�jc��ⷊ�����d����s�tuuݡ.my3�b�D��Nm�Z8�Y����}5+��x�;6q��q�|L���(�+Wg����+�/q��p��d�}�鐥�a��p��Q���WT�����*}~�i$f����)�J�8X�DҦ��mu�[�{1x5�$�y'6���{y��V������&�H��I��u[�=r+_����wfn�4��4�&��v��S��H|"��bf�l�b��9c���-��0�����÷T#�>�[�ʯv�6��亁�Hω�S1߽w���]}b����B��8�X&M�JG;2��5���c��������q��h�g�I����>6�j�fէ&\ �A>g%�O�R��>p�ǸV�HY�`����̶'̣��;��0p�#;׊�B���{;�X��f�E:�ٽ_v��ǩ�̃�M��_�yR̀1v��x>ܶ%�J�I �G��I��ۙR���N��.�"؏��h��ef��>Q���$�l.o�\`�3ٟE�|+K�nY@~ǚ��}��=;�����>�$�8H��.����~	'��ej���Xj>��~����x��{�\��;@�^�k���=�7��T����.�p��3M���N|�AR��LT\�54�
s�]�C��e���(+��%4�F���m��:|�(���Ѻ��;����n�����ϒ��4��|%�)������ϼ>�:.�h�㺲�ZͰs��3�j��������{��b��P�Зb�u�Ibo\F��(Ip���󺺄jv,*z"H᯽:�x�&��W���mB�EU�;����ݛ�"�SǦ�7K^��Cm��zw���Nx��Q��03lp��$��G[�1zn^VH�=���[F)�n�`q����qG�9������w_������c�n�v%��N4��Þ���w�3*9[�Gj�G�_���i����ι=�Q��5#��`ăe�}_q���� 7f�/�w<������k�r���>cC3�t�9���9�o��u���bϢ�1V]ahl�3�i3s9��N~�����){=�(⡮���#�~��*�a��F����M�G���Xt�Ø3�|�ǌzG�r�9X�͑��CN�܌�~�R	#�	R�xT�'@j�	������V��Չ���%�H���{ͥDB��8ߔ�1O���_~UZa�&��z���x�x
N��H��%���ܑ'���D(u{�b5�LV�a�����s��B٘E_�*]p.c�Ŗ�y��כr� %���]�<l�o]%�'��6`s����Z��#=��2A��>�e����L���B��@A5Ab?.Ϯ�2ĺ�b�P[�xs+'��R����MoIi�E�ͭ�C�/�'��@��		
��转��{z�P�o��,&l�;��W�s��0��-�3+II�A�L�H�����p+����"Y��]�����˙�q�T��h�.�>�{��F��������"�kk$�L[���$����>(�h4���gI�{ĝ�ȭrjh���ԡ�\
  �d%fbq�*���0VF}g�� q��J��n��I5X�o�&o�QC�A�0e����:����-pv�X4�uN�/l��� !�׃[�V��4G�R�g��r|��܅u���2�����Ȣc~�+`�牀P��_̉���WӞO��%���xe%ά{bV�X"F��&��%�wS�s��Ɔ����{�����pb��!��W�]'��}1�%Ѓ'�&aDBE�'��_�B�d�58�=��W|�M�G���0������x6���FHO����I�pUf�j�6�r��l,�Zq.���o	�X�y}��4��Xe5
i(A�A.f���$�Wbزm�[�J�ʤB��K��=��xȃ��w��;%!8]��qT������❯f��.�g}\��7�b��)w�4�^�}ї�>lh�
��R	V&�T �w�'gm&�4��Er�]�����ڻ��r�dh�f��D��a�y��uJ(<��z�Ո맶ȋM%#F�����xĨ܊��i����t��UB�� A����9�#���9���l	>��{h�����>��r�a���v���	g��� gg�{�/NS!oǇ�*��qY�$,݇,Hg!��U6)�kJD�na
%!W��C\wH>��ca�?��Nǂ���kz��� Ph9F��S^������c2�<y���(�-zm��q�6+O��Z�y{
]��G�j
�jD��'�ά�5~-�J'2�%2;�SQL��y*�.#��p��)qH��� ��bK�B޼g�\k�a@i .b�,�0�Nt�(�s��Dj� b(L��T�ʖ��y50����t��}#"��]�������1Vi?���4���D|rn�-��X�]FԊpE�x'ki3ڀ�fh�C�����(�W�埣��x۳�w�Ӄ:_��bC��sÁ����oRY��	)�4N�t��X-r�>ن���fP4[����E�Q����H}�7�&Xު�)��!�:k��,��KC�,�Hu	/����򀀌&� ��a�M��SY|m��y�ƮT����w�� �}J^�R�����Y����1�fΔI��K����M��œ}��d�.����ӫ��@,��Q֗�_C���b��w�a�o#siJ�i͂���S��'6h�ⱳ g7)���p�&/ ���`s
��<܎0w��c�p0h�h�5Qi_/̸�.N�v>��l��M�Y�1	�Q��u�/U�*���� �7ak�!x��E�wB\Ȅ���$TB�-?�8c�z=����ZD���B���A�+
~�Ϋ���`���
)�3'p�:�k����N��bݗ��u��}����KN:'Q� [��I��k۴�
�u������E|)Z��y+������"���W�q���6jl�7��=s�^H�ڠ#�r�T����B�{���:���H�z6tn���ED<dB�X����}ܹ���y���ku�bSP��.rE��_Z^5�G�x�̰��W	2����6i^!	�)[�(/�Ѹ���� t�t7�'�>��zIX��y5�[�uW��"��Wn��屁cw�C7�Q�7�%�~�������������� nA��g'�0�1�h�mS��3۷���.�A�N2l�՚�Fl��@f͎�W����8�u׺��q�f@��%�:���x\���d*}�o"�������SL���u��:9�­��:NL*C���ڮ;/������������[����B^����a�5�R	�.?���o|��^��b�$���h�m`a�*��H����PpX���ۦ�g���/�m���b<h(���B(�؆2x�輹^s<��u�'���ow)Tc2���;� ���I�y����K$��yEz��(�qY�5�11�oH�:�M��j�B��7�:�^��k+�g#ˇ)��,�b�Ȋ]��v�,~T�3��<��~��r�w���F\;��﫟�ܝ�1���!̫�S�J '���N��NO@��mZ�q��%r<�Oq(�&���fki<qdV�3�$C�V���5Ig���Y���Zu[�	ў���®rZ�wm���^�xe�����U�Ó�7��ԁn�)k�ѱ^؊y�vm�^1��)V\X��Es����)x�
RNcu7*��u����ő�'43I��b�ם2�}F��2W�y��@<�ic����>N��f�2Y]��Cz>B9��jP���bW�8��- H�D�
V��VS��G�[���~��s�/�����&�^��[�鈘���2��=�� Y_q��DY�Y���G6��Y���QM��9�(����'��9�xf/U� u�.�Rdk��m��k�R��,D&(���]�� H�[��s�
���O�__ �o����
�jxQ.��n�\��]z�s�@5�]t��ۉ����=�B�{���g5+:�<+�[�g�Z/���o�t�T��O�	S��Sǆ������j~K��G�W&[�.��q��#�^�ǩ|��OA�5�� �[G7�&�t�#�yW���Q"�/��{�0�龖���JS|d@F����4a%��|������zzA|q*D5wat{}~��?OωjA���-2h��6�� #�ɖ�׿��s�H��_�ϗ�g�B���/H�F�>'�I���$�i�@���7f�@��jED�~���"��1�qLX� ��R����~��<�7Wb�+� ٬u*��FLC)�?����r�� ���	E��x9��>�;f���a�\m?�$�a)����V�|�Ġ�C�/!��pC����X�B ��E�"��JQ>F��f3 ��cu�p%+~�2|p7`�J�ߜ��~a~�l��;�R�ul���6���	�{�D��[���|��-�Ue�rBAB�A����0خ�K1s��4$ ����@{�?= ��NŃ��~�'߃`���qa#X/tTJ��1aP*�JA�+b�m� B�	Tʪ��>O�[��_��S�<�b�Z������c�m��::���B�}`�ً�.1Pc�V��jd�b���$��|E� 1ټ]��J4ɺ�<4]�ܺ�	@
���@d�7�t�v�����^?O��tR�����ܔ��t����� 9Sxk*[h�����@6�ȣ%k�F���t���O����f�C#H��kSx6�����ܦ\�D�O�Ɲ�a��[�K^�D ��1$8��N��9�GZ�O��)��X�Y<b�V�ύz5�:�gb.j4�h�`�����`�d��"e�ɣX�7?�Y�D$A�CC�viN�2�n{B8�l����f��4���E*	h=���qQ�Z.�� �!'�w�/���F����~�Np���m�������"��w�_����╳*��*v�|=o_�=F#����0�a
8�4����i�K�é�1e^�4`�KxLj�so��K��J�ߖ��.���JǨ`�

��^fA�������7���-`�$� k�/�'�)�P� �bG��,��v-K��ϵ=ۄ(
o`�1q�GH�]����Gݔ�7�i˛\��
�
���GvE�s!jB����֤�v��ω�&�CL1�QH�F�_,d��e�΢�B���L�Kn�~ɐ��n�%��ZO	�9�)��]�S��r�J�n,E�J�@!�EI��	�h��K&�ԈY[^j7�ݛ��!��,s�4Qt3M�U*��:	�>dt��_��&����$-����셼2ߙK6i��6qk�h����\��_2n�Z3�<��+����'�Gh�����q���m�5)ȸv%y��$�Y�/-*�>��r;���N�K��zc�:�@Ǌg��&��ّ?ު�����7�f�*�fjܳ����y�璡�􏑙)!��h��l�AD2���k�w�&����1�/�P��aCd�� �@���<aG��	��?�9��B��>�ܢ�Ã[��a�9(�,���:P��9@��	��p�|�z͊76�҈$PD��>�B\�2:�w�ȵ��K���G�۞�!���_i5wRYԣ�m ŭ����o�B_l�5]�Ԑ� �&��m��3=�!VZ�cE�����ѓ�b�B�Y���${]#�w���"�e����F
K���JVPƺݴ2�an�J���1|ac
��0Y�H�H�����d�qx[%T5G�� sX[��[�*�(�hi��k[�;D�as��m�
M�j����?'��a"(�@�mTҘQ<�.��<;f4�g'?B������	'X	��!��Q� �4&�)(�O����٘c���!��*eJ�%��dkt#Y4}6�H+-qҺ��f��Ǟ~K4Uq0:���=�GrZ&C\Ȯ���K����u8	Zˮ���m�I�IU0$�N�^>\��aYrd��"6F���[�����9����ԛD{˟н�KcX���~�D��78{;�3�Q�&3_��0�w��cS�Q�Ĩ$^H�!�s0��%<�K����
�j.5���c�'����+��~����g�W*��o��,Eyq�@B����/�_I�Ӫ�i�g��c�����?l#ϐ&͈��뜕5fN���M�\�t;��z�E�ZrQ$�� *�؁�e��(�#�l�,Y��z��=^��4y�����3д�%�ޏE���8�"�I%6��}VQ�9�'_xh�� yD�Լ��O������d%<�:��Ơ�~��ď""u��X���*������>�DYW�GN�$
f����	�ec���;.v'��㺽����D��Р�A/t�W��&�M�#@�"R4FN����2�0�ra�p�j���Ѳ�I��0ʺ> k�;[ք��+0r�FT%(�v�-���;�q�AQ�� �!+�8*�"�6yj��:1&�K�,Bpq���J�FBM�o���δo���@p�1��i���<���DSB|L��8LR"�ABw��~]�J�vh��r�,�խ'���G�QQ��Y�%P�
����k��1��Z��"Q	�Nz>�.q���3FJ
ja2���B�(ѣ�=�$��s�0`di��pm���2��+����Y����2s�J˓vmH����U�aRR0L�Ӑ�Z;<}*�����^�ƍ�1�Uо��J�c�2H����F�Qc�|��} *~�P	%��Kt"5�+��I?�(�SP�0|�]q�>2j���&�|�!.w�� T
��B׷ �Ȅ	�S����"1�9����,3��{��>��	� �S��Mi�1�� L���7��5)P[M���9Gy�a{�B��¬Jh��Sy~�8+�͉-����>�@�!a�7#��[�0w�(��O%+�h<�)ƹ��ɠ2�mO�����v�(#��ݘ�?0m�+��|2c�dpt�y)�&�!H,�s �7@�hbz�¤��t�BF/Ch��F��po�����K�.o͎��I�_��p�BE4Nq���q������A9m?���H3����l��?%r��o�*J+N�*J�{�O�8��R�Z6�"	��͢�$G����d���+�kg�
\�
L�n���Fx`xt��+��ݯ�~��u�N>�.3hm�)�CY�M>O�]^�> ��r�)@�;,͗X�2ǡ*�Ƴ˸����rf
�&襳ן�����%+�˞�:k� �4�y����Z;�b�Ve�����sT���Ul��D�<E֑��M��1�_[[{\.��Y�'v�$
a,h�5#��5!�{q�dn�{c:�]V���i�|3�(AE�R9X6��ƀ��"Θ��6 -W�D�����%Խ�ݭ
�W��ȡD�"���KA����[�K����U#�/Ն��+��^��re���#d���ö�m��2����4�_6��_���
��Yp�{���	<��������Q�p3��������qF���9� ��k�:���y%�J��#`�:( l�'p��R��P���<��^�M��UK-t8d��C�����_DO�6�5-2!k�����p��0)5R�y�M|�hCu/Z��R��0*Gv���H�ly	C�3z�b��A	o�<�a� G�:�u�b��]��P`^��񋅚��%5G�9��?,� ��tD���mb|QvN�&J�p���:�5��I]Y:`�8�;�O��w_.�p/o�h;�:x�*s�U�^G�l�p���I<dd�?+���Z�x�mG}���;\۹����v�X>�׾/�k����@0��6F�m��g�/��u�mϼ����Ȳٲd�{�R��;�Y�@�M�$[�~� )
�<:,�d�d�<����^̀T�$�"��{�,D�,<�ijv���(cRm��3Ε5�H�fƔ�L��O8'����Z���S��rc�E�ͷ]��H5ܴj����F�mMހ+�Q���23�5�������'ohʆ�RP�6(�E	gB��B���M�s 4qH�T�`�D0`L�>	�
��IG B~���Qc�!@�v7 �
����!vb���_X��:M��w�����Z�4c��/QM�Wj =��ư�jA9U_f�@9Cy���I+���P`����|hc>(I$��Yoo�΀�l�x���I4� �싸a'~ȝ��'C$)<�Vѓ��%3W)^�i��b:�O��_i6���)���}p�Ņ|R���
oX��-���ޚgH��� ��pE�J��D�Y�@p�ƕ)�Q�XENl�h����rH�`k�5bR��9-E� Ր C2�8������/X�C��]L�
�PqF餝���k9ׁ{{��>Xα?{�׼��N��$>��� �Uz�+㯞b��Z���#+��]c�ˆ[�2��y��?;]����=4��ǯ���lIcS���?u�y���{��)x��S9F��ո�	���,9�^���`M�
 4_G�DLݴb�Ǌ�>�B�ۄ-GfyۇZQX�!J�B�Br��~�$�TF'�e��<\�p�T�7�<��%�y����0��J�tz�$��
�+?S/*x�f��ş�%�b�8CZz��;\:/7�Ql���]�X��l<��0��;q1��@X���f��Ƅy���X�f��1�'k���yXBm�6Qi+����#�Z�
���T������\Ï�~�8�*Ĉ�<���K�s���.̟vI��l���2=D���
Ka���V/�4�*/C�SgoT����7Q�C�]�;�ø��l�o�~*Xf�	�G�/���=�:��7��R�o��a�Q:��mc�x��f�'֪ż�����3H��Cu0��l�J��~9��A0�M���t�$z3�gG�P�(�� �ܻ�^��`:G���nژ7+k4���L��	�b{KT�j�F�� ,������ߥ	˫u%��Cy����:��Ǎ��'�c���c9eS.���	�?D����@�8X)(��R�,Ov��N���f�<0��
e�������F"�z{��Yp�>�F�H�������:b��5^�u�S����1.��!ڢ��G!a�9�B���N��A���j��&s��p�kM��X%x2K�ӯb*��W]P�c���d�� 3+��ε���u��8`��ວx[����b`�!DHQ�,=(����j+�6��������/o4���btF[�6�dm��
?9B >i#��;����|�psם�<~��Y�t��C�A�=B�o��/	j^�I��j�yN@�
zr�$U]���{�a���Rm���h�6���^�wϥ#�]�ؾ���@{=�=:$AA�q�'���(s��W�u�%8ǽD�1{��_�fl��9I��҈"�M�����jъ��6�p���{ n�[��h1"�z��$���67q�AU2\=m��(��,\q�����r�e���ܸ`]�-i+	�9u5$p�^'��9Ӣ�������ӡm��F�6t����v-���o�_�惇�����\�u@������m�D����W[�"�yد���{B��$�������mO%��l7�VW����BG"E�ΨCv{�h`Q���4_��wx����w����]�0�Ed�����M�oS[�%.j,�\.V=�8tz޷��k���*/����m3 8!��a` �xrN%n>�������R2�d"=�L}:ZGV� ��I�+����|�1S���O� �O��5N�|���r+tnFM�U}�:oPR�3Ћi���R���z!^������NWomh�����"D��(ԌKx����Gg�'đ����t�dH�F ��=�������״uk���J}��u6��Gb	ĕ�5���!�j�c���}��䶽[���fΞܭ��S���wG7O�(Θ�^4��m���	W	�ɭB��Cf�	�F���*j��";��ѻ
�������+y���sHF�kśH��xF(�Xh7b�^V?���-c��<Ʋ�9n�9��I��@���YO�1v/<��hQw����)��А�}���;|4>ɜA�������!'C-�9ݺh�7�O��j[�R�Mer�r{T���Φ@�M��Pi� A"'j��֝�f��F��k��I�;0HH-���%���O��*�04G����Ī:C���,E�34����y�.�0���ݦj�N����e8�3ނ��_i�UZ��V����7����A����2+p$)�H��v�S�����{�̸�[�U^w���^��yN�"e�m�áM�밦T�	� ������J��������pf�p|:�W9>�-�6��4n`�L �ޭ�$����'�1�L�)�8�un0Xނ�2Icⅱ���xLA���YA�zش���`�Ҹ-���߲���u�CV��SYcJ�����/h[�v|�n�4�1i2J��*��"/]�y�'<�qQb���ٵ�ZT�@M��G���&�}΍<7�sW���5M����']��{�>�U�E����n[�^j-��t��o�v�ww蔕X�\��_h�]�L�vⲾ�t�;�~,C|��b��=�qb��h̾�2&%�HD��9Lgc7A��Ch2�f�c?ݪ����dԸ�}�Fʄ��*A}��wIO�c��-Ěf�8�o�3I)��ʎ�(]��?o�5��+�~K[�Cx ���!n�h#^=Gu�����>s�n��I晃7`�!�]�$�{� Q��{���s�����t]=��A�P��?wZ�v:p��^نn,�����'���=����f��e��_/���#�F����^�C{!��6�6�۸%�^<n�l��aTv8��F!����}x�hva,��ЦZv�0�����ZK�*V���{&q��=k�b�?z<�����Yo��E�.��n�5��C �wwwwwwww��	�Npw�[~���{U�j�jwg����{�=�g��?�M��(0yK�1�Lv��*u��E6h��MuT�7�*Ȯ�|ȕ�Dl\�G���.w2���-S�q� ~Z����|Lgs��n�ŷ�:k/��G�{�6�	m݃�Kqs��K��I����$�O�l!�B#-��ă�j�y�bP_�a��.��K,��d/l�2��6�9�Qa�㉜��U���/h����l@�%�=*ZK��1W��V�ċ��2�����xE|5��<���)�-�\���=1��}���M�9���k�c���E)�7�V�U����N�9��Ӻ�_�l}H14�5�7�MU�=�8m� -�T�\�J�R�-tA�^�\-��%��..�/i$k�7[-��<�Q�
=�2G�8�����+�>�?�{|��(_l��xU�辆LR���W�����T���@�׏�X��0^��lg.x�����o[jp%uH��!��x$�S��1z�p>��ce�ٌ�k�`�B[r�8��Ka�6kFuD�����.��
e�*E˟TK�#l�D�[����R��Ƒr.� ��Qbv��*Q��P~@��>�d#��yj�~a!7���&�wܵ"�q�m�ڮ:Hg������N���m��'l��V���G#��%dR�呈�㠟�b8��`�̠�Z������Έ�9q�ݎeJX�Q�&�u����au�#t �>�P�ݫ�G�����ި�Hu�N��܄�]<�X�ӄ#�d�ڋ�����o�yL1�S�@Q`r=�3;,rH8!�� 8�,�ُ5�٬��}S���4�,u��^�]A%��<�x�캺N��x_���V����~S3�=X4�`�j{����'sm����m_1��H�UB��Բ]v)Q"��6���3rLr_��p[��p��������BK!�&�K�����wخ�Ko�ٜ���FW��(���"�b�s5�-֢�S��pc����r�r.���ɯzX�2���#��j��d���M#���"H�#��U�Fh�H�ZkJ�_��ߐ��c?�Q�;M��=�y����>"D>�y�� Q:J&�F�y`o uf�L������~>�~��Q 0����͎�_�+����bP�C6JI����T�q���n����u��q�m��j/�?��l5��	��H���a�z�)�q�Rf���iR/j1b�#��/�ׯ����C!��f}��4'��亵;���^d�/��%�X),8,����Z{f��IL���)�����Y���.r��[o�����>'1'&�0y�>���ꕍS<,���?�B�VyJXIe����U�`%69K���t���b�PluUsD�����	1!:���I��� ����_s�;m�3q���X��,"T_�.->`��^�v'���.��Vq������y@��y�0B�e%�A���X45&����iV~�g^R��WZ���t8),��$Ðӷ0ҽo~D�6"�����O�-q7LƓl�;��?f�c�ٝ�[]��[U%�W%y��U�� ��<{�V�ǣ�/J�!���.���|#����kp�rON�}��"3U�#�Ms���|�G�r%��\���	���Y����^P�G�%���y�|Ք/v_:��im���{�iV4].vZ˒_���yc�
�D�Zz3e�`�vY"�bʣ��9JB�E�<�H^�F��k����F��)�@E��]jf��(�+��58�'��'g�R��������Wヂ��?Fz.X-C���N�O�f�h�X��H��DS�y>��hbv?��8��2���g�i�o���)ے{�B5���ds�8 ���)�8b�\�U��|��a�J��7#\�I���C�1.@ߗi�M�뾬A�Y�׉�$�d˟�zܪ�Hߦ
EJ�rIa��J���b䎦�J��a �F��Z�ʪ�-�)d��5�(�W��JQ�P�͆���uC"���G!���{��E�f ��� v���X����і��8vU�m�u�Ʉ�󴡜�)���ΰ�Fm{BC��ܿ�e�?��%bSa���;��;r�ГqU8�� �2Վq$i%��qj0�<�@-5!��}��!�H��U,ۛ#�A�/ʛ�n1=.*����]��.�R�ٕ��H�v�@��b���#��� �����'v �%PCLk":O.�_�7!M�p
�(�h�s*��eH����p��Xi���D� �(�h��E������[R��=c���%�oPzb���b�9�K��L�d�-=�^����b��@E���T�ͨ������K������24�M��
-ǝ�,����o�B�.y�Kvv��8F!I���;�1���{��q�.�+��z��oBZg~���*\�ď��V�76�X3���#�צ�[���Y)+��"�Y�(̎����_�Q�u.��Q�b�:59�jM:f���#����0�����J_*
�xK� �$�`Ie�Qq����yV���f�"�#�0�b�#X���_���n���y�k�O��	�v]�V-��j�S�rf3`��R�ԚY �耱��BN\FR�D@ӎV��]V������ËVR�+�Wa#�Z�W�����v�
�g�3�Mi��%e�'� ��Pm��M���ۥ��������F�I_pI��~�evX�4x���I�ƾ��oK<�F8��Ҵ���������~�feb�
�0�s�I�Q"�}�x����e��T�'�wZ���~,����u��l}oh�>v��������2�bñ�G��{�acMu����ULw*z%l��bsd��� s4��7���ƥ�q�ُ�&�[{���^%-����������^��s�n/���.�$��b��%lG�?)sOh�*4�M|�N��#�KXJ\�8X�0��5��Ѕ=�{�]���"��nfJ4��� ��L�(��#D��9Hug���@(���jׯ녔�#q��v��HhM9n`i�����n����Oi�n�w��'ʛa�}3n��N" M(��3��6�L� =�P��9���n��n{�?�7�Ȓ�e�C���c���i���E:b���)�[�m[qVE�����cjd7�G4��?g�v����u��g�E�ƔV�A���>0���oT�=�_��|bc��@���&�ѹÍ)"N������7S�n:�;��M�ͯ�mndpWt�h���]f]�����
2�?W�^g��øT1V��τj��;��Hn
��Z�P�&��ݦ3�p�8��t2�5��M�haޅu�Rj��5Hy���.��^������h/��Q<�<��\�ԓ�D~�La�N�F�� �������vmK%����-mȞ�ŷ����8��^��GN�2ρO�2wV�O�4�qFH!]^�
@�83�@)�G8��8�K�9�̦��s�ӓc,�_h
Y&���P�=L���um�ZQ�lo79��|I�||!�QZ�T�9�,4�5јVl|��T�y&I=��|1k�%�ل0S�"c��~�+Ľ����|]@��+�N�ã�~�ӄh'����	{/�.���|tĎ<zJ��J�m^�R=���e�Q���z�fg�Bգ�:l���X@-��JP�t.�*>�8�����}��K�D�0�,m_��"����l ���9?|�'�9)�%.R?���˙�W0�P2 cb�%�dm0b��9�l���O��@�,L��%4Ɏ���J����\7�E�=(`v���lP��Wu�2�S�Y�Ğ�lֵ�8���:x�z������*��S<� ڱ��agb���Jv8��s��4��Q���6?"d].���F�����С�|�[�)��H ����r�����2D�>�FѰ���KU^��I��h_QRE�9oO��8:o�*l��ͭ�-.�w���9c@����RL,��.d��$h��J�X�na8�1�Z�9v0�^ى�?�T�;F[jc�l�i0q	��(4�3����ߣӸ}�J�y1>���W��.�����	�#^�����똉J5����&�4`���~�e<@[5PE:�	�^ǫ�~ŕ�c�?E���p'T����_Z�t�@��5(e�٬��JW�1pg���%�G�}h�-U�X���af��q�b���<�-���[�=$�
�,�����+��+�a��q��ޏ�g�;	�;&��d�_p�4tx���F���2ܘ]ʫL����}�wN�<Ԋ�]t6[y��Ȑ��9R>`�����7��H�d-����T6TǀҾ`�&�����|UKsy�7}�I�7����Y|5�{��9a�x�p���*ineu���׶1������#jT�������*~7~j���t>I���� Q��j���7��ō9J�u>"D
͇����0��� W����[*��߈B�+ ΢�hDx|��h�b/ڑH:�� �nCC( ]���8_A:sGH���q���X���l�Xo�����n�&�m��iL��ٺ1��'-"`.,�c!���D�w�����J�����D��ZE���(��N�*��Ǡ�,)GE��}��{/@�/x�\u��,-b�0�G��_�+�%��]�\7��a,<��e\�-�n����խ���o@�����J�滋H�"�	JD�M2��s��Jx��t�а�]�����$a����-֚R2ʲ��Ώm��i���-p�Y����O��24k���T)�5�U��L�^��-����E[/�W�&��T~�xI]�p7)Y�GBѲ(�o��)�I���^;U�[<��7���P�V?�Ŋ��%�i&�թ���Q��L[��d'���؜|�3�&�=�*�XMp�?;J�Mz�x�m�2��(cuz�جG#�@��f�R�\�%�қ+���-!��[��0�֎�y=y�j�=����>�;y|�v+���-v��{i9���j(�v9Trs�->v���V��q$�\���l�s1����IǇv��0s+�ϮW��S��R^�(Ix��L��m~㟹�%Ć�q�GH'�|0�6O�.��>�e%w
f2�*��K�X*��̮D,Q}��~V�5�����'��2TR���v!J��w�������7:�'=!e^�>^!}|�{�9W����JMa?nJS���P���1�l�s����wKo��UZG�G�=����\[l.-�7��M�q�e�xjj�o� �CiV҄<7�����ќ�K�,Z4K��K�ݶ���ވ�:Z�oNbS�^��#��-[q"�N<i�!b�UQ$���\c�۟�Cs�W!x(��G��U�)a2v��5�cԊ�c�6�I� O9�\�]�QEk��2'.�|��u��wP6a$ƅ8�EH�|^�f���_�g'���ie-��FTWĶ�_��Q��Ir;#�;1�~{A�6)H��%���/�bb9Iϙc�W��1_m*W0��a�&��t��S����Ҭ.C�6��)��oQ��+`�CDp�Np�c��̘�3�tI�gO\}�����q�{��l�]V����%sb��t04�X,
�&�,��ف�/&�i��e �f\�1"sЖ�Z��*l��-[��[�a���E���:�] gr'P��7":VD����?'��;c7<?�k��H�z����iP�J�(u+w.�5�w�6|���@��S_]���	�~�^�o���Ϛv#�kxk������%��A���ҳ�X�ɉ�kK�uGE0�U��~ǧIߚk�tU경����hh�l�a���B��sM�s�rp�e����� ����	D6�;|�yt�l�X��9�ǃ�dT��H1
Tk���F��m��	#{b�#�E9L�a���'����D�:��S,9קϱv�$K�|�V�q !�J�sN��S��%aD)!� B$-�|c�f�'��"x����d�y�\���#Y�����&{�*ӓi���wֆ��\��p	1,��Ѩ~��*n���ЛX�i��[��<ZD��g��iU�-��V�n�Z((Q�A�I�ۦ)i��Sk�N u�F�L�1���
��Tl��i{�|������Y!�;�7)��ӱҳ��4�S�(�+M�Nm-��*��_!�r�z�B�[y�C�2�\��{�#nM�qIv�1	��c����V��b�W�h�&�H-O⤯�3�N����d�PA����+��g���'</������B�P$-�̼�`�[B�0f~O�z�X��;=vKs���k��&�������A֕��*߻�;3�࿺?B�q:���i3��;)@�S�(��쀌�I%҉CE-W/U�����9L�=�'��pY-�����X�uQ$ѩU���E/�DQq�fW�M�m>b���)Jmgs?@��A-�o��
���l�j*�*]>�$eǂlu�ٵ��5�Z�e�n� �"����+{9F!��1g�{�F��
U��`��)�'��%M��#\�sk`�SĮ��}3���1{��&�^�`'y�J^MY��?
$G
�$�'�"b���ha��o�}=W���`�/޸�ӟ<Ae���me�����x$��h	h}m�\�z�;���u�nBCs��9�ޜ�6nU��)8U?�,f݋%���I����Q�8�y$�"i`�^ұ0��뚧^������Wpc�l��5#�&�6B���fղps���qpi�Y��pv���um	�MRF�*P��#�,!��L��GD �	�2�X��e��������o��"�_��J.��Ԓ�d9�I����B!4��qw;����o��ar��($�ĥ���LG��f��UJ�L��E���f�c��,���YrtZڮ_����F��^���B�)pw^�w��}G,:��PC�����m�P�rY�_:�%��*�Tz��e���R1
�R&�c&#�&
Pj7J|�=�,�ӛ����Xy��)3Hb�7d-߽JĹ:�ut��D���4��~��w3��[浻���3�$��bY�ܟ���H*�y���cdKS0~c��@v3��Z��d0p@`g�p�c�#qDSB;����Jk���K������ލĪIO��+�[��M�����E�=5]L�qO�f����v&���,��\&�����&^��"wk_�6/�����'��ݕWh����F�9ոq��qL�+���ܨy�ti���]�ᢐ�ow�2Q�}���t�襏�T�,��ދ"rz���g��{���B�΃�+C�5�,y���k0@0$.
��b�;�laS�M��//�|S]��&V���-�\	�
Ib��Q���"�wg|��x�z���H�w�Υ��;��KiN����������	��-���?���\,�č"j{sS-͝{���һc��q�� �)f��']��-g����(�O ��S/�f$»S,g	������FN���j���u���9W�7� �=hHͤǯ���m�� p�}���`B��W�'����b�t�_>�_�D!�Q����4��νkzI-�L��#�Z~�;)���q�
=��P���%N~R�3J�MU��٦��`q����j�<`
�M&�ȃD���Sk����"q���f���i��tv���s�(0ahG�,����1/�[�����:R�"�-�ʢזk/M�k�߸�ܭ�G�M���+O�3���$�zЕ�{a0�+9E�ύ%B>�~���..�B�%`/:A���M��+O��[5~�[�3��_�����BvOe��e��K"�"m��D⿳甏����5j��g�yƆbu{�����Z�X�=�X$}\�.�SQ-�����/7E���豨5�Y�%g`<�~�y��y��_"�k�P�<�@�p{<�'�m��(�����T��m؈!*6��1�s��U�Gߑ�{�������W�	�qDTf�,�eu�@�f�������R\�{<l�1�<�W}FN@N���D;x��b
���vޘ@#�֞G�s��p%��B�׏�uW7��B�����*�ƭ��KC�zeGТ�Ұ���۩�\�A�E&�)_2C0dKj�3��<��*Mʛ�2ul����gJ&��b���o��֩��:�.x��!rq��:?�+��ä��\̔��ܯvɒN]��Lǝ����9Y  Z1Ls*2�m�)�J�{7�|����~����f#��A}�������nh葅*:<�Q<�g����3��j�v�0�ߞ���_-o������t1��P5fW�Q#08�y�ں�����'�����b%|�dz���-]���A��ҳSgɪ���x��G����]�=��>#�n������z�Y�$�$f2jYؼdTk�j�Ȩۺ�>��H��Y�z}�'cv��S���Cbr�0c]��zb�c�S{}�Jq��R���8s~'�rg���z�_B�_&eϚ(�&����k�Z(�'�L���e�yND��r#sf"!���.9´�#������N�l�W��0�>j*Z̙��l���|$c��.��<	#�K�t�%�]�w�W��d6\���E�!h��cQ���+TǱ��J��)g*�AO#߫)@�F����#j��Dv��8�1�#�������
���������q ���C���{� �Ĝ���mT��N)�bN� � u��T$h�TA��!�O0�>;
m�l=�+9o��i	$ĺ���L�9X��]C���!#��U�Ow`���_��u�1I<B�G'h����j��ȇ����������;�y�/�c��M4����D���Wr-g���TOT��x�Wqɑ��	{O(A��a3�\�to���F�l�d�)`�/���9$�1Sy � mؾ4iYzѼ� 2�N-U ��v
�� ���O���w�G��O:,\��z�|���������=�U��W�K�?^�N�9��&���
̹��D%�.ѐ����-���r/��8��0R�e�����3�t=}98)�PY]tb�1��K�U���&�-F��:YAyg&���'�?_Y�[�C2-;:$K�J)~`�SN��8n���Mi	���%	cA�����
�y���?W�B�e>Uf�t�({�����d_�\ŬI+#+1;��fD6��Y�Vj#��Y�L,Cf��/YCoȃ��P�5�AJď���<a�X�����Ȭ���SN�L��z�1r��&�p�3d.dm�;�e�_z)���?���<�S�嗕�b�/^��A�geM�R$D����1�Ox�!��3�#pKv����aT&;��U�c)޿��8/�����%%�h��|�j�i"��@#����槟�ŭ�
	ꏜ�^{BHaRԸ��r�ɼ�{qq��hF��/r>��~���.��G��f�G���L�LYk1�qY��g�J�LS��u��P�!pL��_{�Ĺ�P�ٵx����nL�n#�z?��q�[/�Z���*�����"�c�����e�]�{�2�ȂPəE0����,5/ϲa��җڌ8U�L��6��W�2eM����pG�3#�5�|X��+���"O#DôZ��5��pk�(�0�e�����0��M&(j�J��䪟�k?�����dْ�ēz����~QT�͇�������P�]R)�;�P.�nν�ϻ.��Τ�{���0v���B����¦�m�a;#��T��=���͗�&+���ݷ���w�8Ʋ�<<מ��41+��+{)��z*~��ASJ2䍄KV���JJ��&m*�9�ЂT
8  U��ͩAEh|�e�Pj>����OW��9�T�}@�\��9,�t40ș�}g~�p�K��*hV�)�$)���>>��DC���E�@�x�gE��1�X��s���i�E��ؔ�6˻�Iv�l&��r�����& ���筇j�k5�Ъ':����-��o�P�g�����c���e:/;Cr<�#'����w�=��H��0�L�hJ�~ ~���Qo�)�Ջ؁����?oMtDx�1���g..�;G�z1�R*>x;�u}�>����歐"ah��[��x%@a����|�������(Ll ���/���1izI�!�4�:(���v0�h�����ï;wU��{�6|���{�Qq׫X�q��Z�m3M��1k������P[p>�����V'hP��(p5��Q���,�� %��+����&eg^��������L�Gw���X\
��)�q��r�O�$Vo�������'�4�7˂e_�ּ�_��2k��-�1"D\�)���
��X���aq+m�(��u+]���G1�*g[�k5W��^�������;X�ͭ\	I�@"d#Z��4��K3��
��Q���U./��Iw�e|z�eSl;\������x�:K���J~Td��>���r�uPuh��ד�_1�#�ƨ����kbJ���p���" ��t�PW���u*�&�I��4���E~z?'Kǉ+_>�߭x�P)R$b<� I�
Il�´]�������p�:�[���������PM9*a;����z�PRD��>�਀����=���p\��v���N^
LxLx,5�����G ?=?1��$SK� �ګ]��*F�l����ϊ����ˡ���]���������~9o!X���Je���-��M40ޑ��D~  �VLPL؊���WH��i�F��hX�O�=�K/ �A�%��Ȫz6^�R��q`0�bd��ۥ��x��b� ��Q���<�ta�N�qX���H<�E�-�t��L������F�J�}�<�0���%�v�8��v<ѩ�"��eZ���@C.O�������`6d�[�� ( .�����F��%��'ؒ����Y��cs�m#EH�/�^G��kik���ʡV�1HmZ2����k�����^9��x1�"�˺�~���V�Um��ڢfG�
�A��(�D�__B]�U��u� X/��������nb̌��H�T�P4�+Ѽɔ
�e����fz�-C�K��WSx�qh�儚��m��0�\#c�&:cZav���ƑL�eX��R�_8�Zk(�(�MŪ��6�#�q-��~�����	��Z���c�MA�y�E3����E�V,[��(s_Sf�ik�2�>��SA����cg���E���ݍIU4������e���\� ��_�Ѡ3��������%S��T<�(A��e�����rG����J����i��[f�v�0:�D�kE2���m�F�B�m�K� K����B�x��x��@�7�g���ŀh �2��πx�`9b�	3$3#!A�xi���Q�f�'�@r%����u�#Z�cƔSH�n�"����#{��O��CVB)=`d��H�U
���d�����&i�����W��F�Hhp���)}�+���B����9J�������Y�>z$�;���IH�(��tc���^ϊ(��k�A�[5��:�b��)������ ��mPI�g!����i�	� Ɓﭡuud7X����Q�Q6l���� &P0D��k�1Q�1�ݠ��#U���/��	W�4�~���|����������#0��]I}���~22�8ZN2��2#q��|�P9	��=
�H/����C]s���O��WD�;��B��f#�ϻy�ʳ�r?\�ӻx�y���&���pX�#���ٮl/�cW�O�?xF�֎�֮l�+I�+ǁ5l�~C��|׆�zX�jF�CՅ���?r�?��$�%��[%�ȋ@�zbB^�L�����(�$��͛ޢݪw�@�:߅��Txa�p�����p�a�XwJ�R�':��!����Sb����P�|h/n�?)�5Cd�,��Mb�ߠ}fŊ,�W���H�|+�0�^�:�;G������Waq�~�_��/4)��E���Ç�Aq��5+Uho33��$lt����S��|qFJ������9����[O�g
T}��8h��Q9�P�/Q!�Z�י,ĥ�߆��A���q��9��cbs��#U�h"���D�5�����季47i�Pf��ry�L��-���y��u�gcN ��R-��<2�����-+�K.
�������m�p48(��bwkw��/E
�b�+�p�tL����,uP�@�G}�LfE�"(ѽ��9dm�7;�s=�bD?�nD��f���6�L~j��n���{�׫᧸�.�uю�`�xΨ���`oE[$�����v�ؓ���r��^�ʙ����<ݩ�1X�ʐۇ�ё1��a��M�r�)��=�7���eOj�_�n�[qVcR���k�"�'RS͆^t�q���6������F5��Ϯ���z�X���f��l���e�f�:�>|<�?��{�|��k
 ]#�a9��F����GBKb+��h��L9��x��K�Cػ�������2�<8Ć��y��u�^�~�7���5q�@w�G�d����;o���oy�K.��1�}X��QTh��Jܲ���j�H�M���7���-$|��\>O]��(���ܽ�7�2;����y�<>(m�w��l�� &��X��V�$�"i�c��	��K�Pt8��5��5���"!s���Aqpb`�}r��;@���Y@����T�P��ϡ�j`[C�_R~�4aG܃���n$�/��������/U����W�߆=%�-�B>O]�����<ޠ0�[�.X$z�`���>�XXx�Do���0����sx��T����zO��f!�/�VoC�QZ'>��5�;��p�����٠3*L���Y�Oɛ�/h=�(b�GHl"0�,x�,�	$o7�AHm��,kM9Tcc'6*�V��Q����LM��u�X���t�p1��x��s���"�Q�k#��� tRI��.5=��D���"*�G���n�ϣ�DC2���WR�k%R9A"��w��

&TM�0���kZ�g�#Cm0<ZJ9�䢳�j� �:1����;���n��GJ톌�hS�	A��/�(i!Ԭj
Ʒ�XQ�n��y������\	�"rҐ�����U�l�@@�耔?�U���$�����?뚌K��,��7��#�<Ba�M���c�������	v�j��Bl�����������v%5<b=r�j����ك��3�Ա@�b������inQ"a#נ�a�$��.\_8b�n0��ē��+� ����"�Y&�
V
�n�x�]`��?-�@-b০ޭ௠�h��s�&Ip�?MP�YU��_�U�>�D�W�'�^[͸��J�7�� �\B�!�����48�9��̥�F�:f	t��vZ�]�o��q�a
������՚ax2����԰n}X���Y��^�A���&5�M�
�X�O=^5��ضN���*W� e�����4u��Ll����F����n�i���h������0[H�]	?G����@.j�Ttàı�+d��rO��� �c�-��OF�+�T��ϣ�9X�
3��Թ6J�軱�i&C�G�Eώݘ��g��I��\J+(�z5l�s¹3q���2S�b����ҹ;\���F5�:oF���&��0��!rWf��5��Ħ+J3� "�{��P���r�|�Ⱥ��B���yz��%���LF���o�`��M�T͢DE�zp%�
x��[~����$��i\f��1�ǖ!B+!|��_�(-��.a�O�~҂I'��Q+gWF[�ȉ8h���~��{��;-���9=ul���W��N�v+�>�z���*�R9AZ�=��x�'����*{�[��k�䷴�� �bu!sZUC-�a��g:p�:�+T������=�Q�v�B��@�S�t��R�ڄF��^橜�e(��݂)��1�����t׮qiΟUmڷX���=�Nz�$H�9t���1X�B�X>�P}�?��d\��	ʎy��xZA���1M�%��U)�ک�[�U섎�@gB�Y(d�7}�����[Hn��lPQ��2vvĘx��&�i��{+�X�"�'�����=2
�i�`�U,b�gf����G�l��"�#����xI�;��鈸��A�,5;@F����*�P�m��&���������V�k~��K�- ��p���x�n:�>t)� x��M3�)�M�l8�-����KG����8�`UI?���`s�F�p�2�}Z�����O�Kc�f�
�!pӪD%���׷�H�
�8}�Q/�`��>z;C���49fjEPo���X�Dr��;�5���^�[� A67�>X�R�ny�7i<��PI˞S��xMx��n�X�_��O4�d׽�0[Pr�eT��⽬�k3<nvGV�P�^.�/{5^�r[f̉�6�y��y��E�YE�G���*���Ur��%���`��Y
�Ʃ�@�����F1n5�}�z]��<.�W��D,J�d銛a݇�Toud���:D��Y�$��6�+i*$�C��`�S�ws�c'�]!L����qZ0<��Ȃ�u�Nw<�����D��Uo9�i��ş"R�!��,;�6�\(Ճ>�X�>�"\祫=�Ǿ2���`����_i��S̹�1� :#��j\�����[�'��f���ن�V㴴"veў135=���	����ɧ��� M��`���c�5|J��i���'E�)27�J�㯐$b�)��B&)U!���f��A�m�4�!b͆�qi��}�����J��9O���n�8��
�tF^PG���x�\�x�[c�v�RP"?SJы"��q�r����$��Y�l�(�-�P�J1��^	CM}h�T0��	�P�Cj]�P���C}a&��l���Rگh�����@H�.ޮ<ֹuSC�˻Y��h�Ш��R���.���=�C�X�;�J%V�ik�W���z�m�z1$ވФF^�7^�'ۂ�1����j�B�tJ`q~g!t )c!�B��|�-�k!�Q��O\�'��72L+�|��[9�VX�7ڤ]<e?K/��@/W�Z ���d_-Du?Z�s�S2�&:�#�$������tJCe��U��M��;��F��x�jdwv��ѐ�8��7�
�����1��9�-����"ɅR���48k�nն-��\d�p�=��zd)�hk����ۧ��+ �mT�v>�w�t��7=z�ʁ� H3���F�K�#L����@l�[Q�����6�2d<���'D�T�F���-mV+�#�&��0K�R���k	׬��P[f�_AnWL�ˑ�U*�u����$�zfz��F�Ah���B�Ǌ7x����ݰ"�ne��u5�B<7�++�����20ŎW�6�<����ܑuk�����\�@�B�)+���k���M���J�\KFg�"T�"�E� h%�#�T�  ����x�B�,\�b(g;���}]�@~ݍa��V���$��]�+9��FM.I���7��3Lp�e��sfn϶���bs�+������X�4�y��� ������8�����"�$�	f��ri�3������MǗ�W*����P��'R�t"V>�!H��.�҃e��8���ܳs1�� �뚋��k�6'}b̧���3�!.ko/DK�[Q#g7��e�
�E	�zzh~�p��7LP���-fv4��?�L������5��zw������Lӂv�~�F�:xe�~��;R�r��|<7Dת.c�~(r�h�r.� 1O�$� 3u�fj����(3m����N�>�l�|o�)]!�K�r��?�F�ڋM�~��u�������K�$��8A���F�ۂB����E����z���%:|���Tcnt�Ve��=�)[�p(���O>2�W���u�m��Nt�>>H����_C
�k�S������I�/��l�4B(������Q�lcNx���#S6A�s�d�m��6j�-�-,�C�7�Mr�x�61/x ��QPR�L�㱥��;�m��(=���
�#���ǥ%Q>���/|��O�,����F����\T��L���k~j���@�����u�.�"	������G���Qͭ��a��:��e���>�6���m�NU�1���a/�����d�-�p�ȟ�t$*x�hgl���{X��[7#�3K�*�~��Y��RN�7*+�	���J����L�������Ȏ�rO>x"�.[M_�	_���/��SD3���/�K�+Q)�РK]���ճʈ� S�K�gf�܀+�D�k�y8x���o@ݬ�	(����|�#� w�8
l>��������3
���f&����Z)�ϲ�"a��V�����' �=��e c�8����]������0�O�h��y�"�������W3M�A��\0)k�ET3�q�0���>ҳ�=FY~>�����:9�_t] �;�ne��O��/�X��R: ����uЛ�Б��ۨ
��na��y�&�{�RO�]��p�>��[
�R>�����I�d:�H�N�1�ż��՚ghM��h��_""���<��lHaoh�/RW�;%��Q���g�J�r�
�F6�1�9x�m�����+���0ww	��������5��;!�����n�/�n�{ﮮj�v�gG���z��y�?(訩P]�Se�[�P�x����8�>��R
e��c^MI��T���7�#�ʌt4���h�#U��NKv%�9L�U�.��9�U����6��V�B\�ِ��H��b��}����"y)��tϢ����m�[��^L~ng�p���;D��|�fYg�՚�Z; -<O2.���{�;�� >���Sr�$f�X�db�ߧ��sP4�AF(8EH�v�ӧ�%��&T*T�u㋐R�tI�=�����U�|L�f��]xL�.mL){Bh���$�-)�{���ǩ�M�++�M��d��G��ik����@%߬5B���Tk��#l��$
y��f� �����*~�~	�h�*=Y��fܢٴg���ǐy�Cذ�	gT�F������~*gC 54�C�/��$6���y3�^yG���>L��C_���W#2�#���8"�V����z��hm&7��sD����T� �e��Js�@��OC�ov�$t�)� ��*�@�Xտ�$�����%�Ù	`<g,Ql,�����S�2h�U�|���e��Z2]C;���s��N�7ҕc�~�Q:B�$C[���F�dn@L����X��/��;i����%��~l�*���L�G����k�
ޕ�F'�)�1cD�9'Ș���f$���F��ؤ�W�_�c�>oz�$񾅴�E��0�����*�7Su���G�]��3(�U
��'�@x�*-�^чY�ʎg�!�Rѹ|gCĞ8�̈ޣA�
����o�J�%�)~�R�x�%I/��̷�I1C<��20�kg��Ӵ�l��i�d��CM�3�_�D�<�|e��O�kII�_%�j�^7���L��ߐ7�T����B�є�D�C�|�`(����e�B��8�-���F�G>��2�E�	���K���C
�t���$C��;�5�uQ�!.rX�W}�҃�YU��8ԳZ�&�{��ږ��x�v�Nɬ�;S@�G�P���%���d���x�|g�}�t�a�OWC!�R���~V+�P����o�HkbX-\5��՘�H4�%e񵓥����~�����/nO�[f9�n���	�,	�x��r��Qgְ	�(�pH��$�5n�>(�}��'7Ϭ�{q~�솳Xı���!�\�����.$h>� X��S;ђ�o�~����a:��c��pzT��榳����\|U0L;���L�pK��%���s��.���v:k6�ٱ�R���T���3���Lsь���K�o�9�����s7�\~�C�f�*�h"m�QQFK1����V�u�0�,�#��Nvc}���xC�9P��C�_8����^�&<`L��E5�ٽ}�޾%�_zJ��dP�7��C�U{s�SP� -�e�l�hG��p�T-�Q��:��tw��d�f��j�\�"L�����'�е�d�з���J�P�B-�Y�Uh~-�� ?nrN\���8�u3�7�z�^jԷ?�_i�uJ�~ū�)�����nL�]����`�:`��|�թ��+�l����+��k��'�R�h.��;���**#�0��,�D���78�)��%F���EV�*����C5@����P]s���	I��Q���o�i!=�A3p�h��I���
e�߰R�y�oR���KF�^R���1�����y���� ۛ�I�(Π�W���8�#m)K����ۃ���x���=-������nS�8��ܟZ�&�D��4{d����;:?d�T��z�����k��I��Z�����an:��ԌP�����7�g�c�fE�5�[���M#G��D�<U�����S��0D��ԁw��+TDi���)6;CF��5y&Fzc	2�sr1R�p&�����鮆R60��T��s��\����|�~��������U��cs�ϝ�>]��ރ=.�i�g	���n�x_���BI�L���IoƔ�C�^������RVDY���ܞ�����5�^�
ˏT�|��5��T
�Ԃ���TTV��t�G�)���6>e�|g���	I8�Fm���S���^[�n2@��ݎ���R/O�+$��nn�-�@,	�����}���`n���4F߅Rw�� |�� ���X%�R~�T%nLO6	��4�df�w��[��,!�[Du��UŬn��!-�����u�N��ςz�m��\9����wh�`i���,�Ҁ[jz�3h�rLJ�0vۄ����[h�+��FE��}A{Rp;����~f<t��	��Qmk�Ty��	����ַ=��AcB�%�#�c�8
��?�m�v�	�N�VT�3��C��}��Yẜ} 
��(J 0�C$�V��+	\�w�%�'T����l<��m��G�#�Y�.#>a�X5��q$��E�����D���`�{+�#,��:yi�8�=)��嬿V޺~��m�������:b�E�$�*�Hۆw�Z)�n��t��� �p�!��q�B�"��椴�X�Bx/Sx#��4x���4������*�ɟ�`@;�$� �zU��M�(rtd
��u}��d��/�J�3Oy��T��s����l>|p*䣆j2E����"p�N$��H\h��F��?֯,ܘ��P���+R��*w�P%��o�I�i,׎��a�ƫ�������$	�����.�RǦ���>���,�D҄&���G��k���w #�
á|�6�µ� |R�._@ _�FV�>>W#/������_B>n�S���J*fk$p���|�K�j(��8�Xǖa�x��q��eG1}�3
�//I�:;��	\����8Zr�����rE/�t!@fu �^������?-�q�I�F��s
[~�����CS,&�����&�0fp���ٯz��H������=o�;��vgUř�WĂh�@�5q޻�0j�d`�O���ձu1����e�y��!��dZ��`~Ÿ����C'�MR�t`��#h�#.G����v����*?/�����^�
�N�^8��O�2������&��6d ��w�m�LK�c����pS��Z�ڨՌ+KP�`p���=�ТY ���1W��9V��?\�����\�R�\�V�s���-��av:}�*�����[�s9����EQ֏>�/�	?��f�̻[��	�!%MW��xm�d"�Q�SJ��� i(�A��~�Oo���#s�&A���|�ЁDϥs0>}��r!�*��D4˗5(W��|��W>�G�ợ4��f4/��e�s��l�I��H���]�t,ymo�~Տ�Nr��t�=�Z`n8�4���k�L��Y����������{vN8?�0�z"�G�W���`<����5���>�,.��(d[3B�:K �;E���`C��hO��,�$�J��"%���X��q��"�.v1���iP���Oc|�C���.�+�m�c��|ٰ`k��ƈ�k$�� tC�e6|nի��4L�'>�t�e�-�$z~���;���+�ֽ��Rm���ZZ�w ���JM`��&�Q��h@�U)%���yj��0�G��n��eo�~��m qE;C�;# ���/���B=�,"�
'@�%��G@{���:�J�:7��E��=���Ly��s�ߏ��\!�~sv����F@"թ���5���"�I�|����n)�&�ϡ���s��9Tb��OPվ�s��"s^�5�%�A����D��p�FY��O���Ѱ2�rI���h>������s���]o�TR�߽�u��z��������t���"��ڱ����?�p�a�fT���=�r�&Y�ݑ!����S�G���bw���k���(o��x
�d<�+&m�D�"�ȰPK�{��p��ѡ��M��S@�q}�=h�ׄ�y>L�����깴u����A*W����0K�M?�/ j��m��{T���>xVf}m���rh���\��\�U��pl�XE.�l�H6�Js_����>������8���iX6 -z�˴��n����MH7b�����7[8��M���K"�`����d is0I�hQ-����,؋�Z�:c�ݛbqk� ��{�|�����e�������M.s�����	��3�ϥ�� 	hW��9с ��k�=�|8����ȡ�X���Ĉ�s��wmQ�&R���[�^t��7��m�%�u>-iӌ��V?�`�����c���ܴ��x���OtZ�@n6ȁ��o���ra$����\|���)���s@����)����/�$�3�*	��f�9��uz��
����n(WG
0Fj}��[@<&���q��lq�L��[{I	�ޝ+���w<�����KK�Ʌʱ�ރ����E�7�ű�&	���%��-lHZ<����t������PX�mݤ�����d$D}K��5�%�+�L����Wk��mG� ���]�)��G������m��n6�L�f��[IX�}T	�]Hl��(S�����:=gư��I��۸�N�'��]�!e�pG=��Iq]����C��bܓ��U�����2����+m��{�`jq�h�FYv��Ajn.|��B�"0^�.�!;�<)��\3ˀ���.Kjr"�gCu�md;]i4m�?!/�ܾ�$��N7�X��1���CDOBM�8k�A�e2-6k��&�{˓��Om��My�ywvv�����H�|�)��TgF%�'��=k��=��ïA�`�KQ�ZT7q\2vk��U[�!��7O?��]"��a�n-��:�#R��������)�x0�3_f��
�D
��a��NoM����wx^���S1� �߲�.9��_��MK�v�aJ�x��d�
�,Y�X�ȫ��N�=�]�7E�3�E�l}J\MCV�#�b�>��=�CM7���c���t��A#/3W
����M0�[VP.�{����9�� ���Ck�O���h������OvEߘ�̷��&�I����E4WcY+���s��.7]>t<N@ J���g�z���Fce���)||�.��Q�5�,��*��$�C�v�Z 範g��d�ໂ�z�-Ԯ�#�a�T,�h�[�*K�P=��C<o����u��B,��	�N�����k��6�z8z�y�L�ʏ��ټ��S��('u������hؓJ�oع�ȅ!ӑ$�O��JM��P��!�Y3��Ƚ�3����ɟ{�,9�{��Z�����������d���:�Rˠ��%�e�bg��uD\𖾇��gf��8���
�[qI��d؜�P�.����4'H��P.�Q%|t?��"�w;��Ҽ5�D�l�&�Sh�J��Q��F��~L?�ȉm�s!�A��Z)�޹E��{ۇ�G���8������{���J�� ���E�#�������Rb+�4`L6�G�|��F�K?��r�g��IWйH^�q-Mn�s=u�۔�d���3�&P)�t����O������x����I�g%~6���Y=������5�9z1>b��O�G�w?Q�|�LP��l��U֢|��#Tc#N:#C�|�v�\>>�Dk�W_7�&P�+����^�>y�ݳ���W'�Dfh@5�³mнVe����[K��B�6���]���u�JJ�B�:9e�q7����/��3*�r���8��B�GjwP�G�U�)��ſ,��:W�;��qaݩ8`�������%WQp�])���Hʼ���G:� ���ViN��S�D+��b�6�?�a���3?]*�r>h��<��������݁nX��"r�*���Ɩ��˕|� Z�A o:�?�x����>2�~���l�#ξ3y(��3�V��� �Ԣ�
���7�Ᏹ̙8��L����徾��q�U�s>�p-�٥{,�˔x��g�Z���]բ���/���,���՝���qsu��`BHþ����5�[�ԅ�������|�A$�a6�$fB���Q���5�x;�F��G���c�B�
��6";ĺ���
��oW/h�3�x�K`����\c�Bם�ul�s�)﫠et���[�U䌄������&�܌n̯g���(`�E��rqqI%ѵ�n��G��$p������Ͷԩ�\ �e���R74990�؂;�+ֺ�����W�3h��էBO;/Jb��<��������[�j���刍3�cM���B���⺫�Z�|�s�7��}�[���Sjf!���sy��`\X�ɾ�~^�k�VeI;5�=R%���V �g�#Tk���C/��i��!KL6����ˤ�h-�)cv�5�g�QB9uz�>�0D4к������U����u�aA�ns�KE���Y-���:P�I];�����@���/t�=.�r�6�ʧlj/}�'_1�
���P��7� ���S�l�����r���$!d��tpXr"�Z]�]��^N�(@���9��t[�Qvz@��fD|���$����Q��{`Ne��k^l���`YJ�=s�%oqg����������៾��;��^s��ȥϴL;�e1L��(�1|��{���w9!n'h��'�]3h�]���
�
:NЋ������|�A��wd�(��T9�c�s��*�M�sd�����7�To�a�.Au���H�gZ <]��ĭqǍ���C+����廁ҷ?�ڪ���&�bp�)~��2�/ʸ��45�e�Ҩe�h����3߹�<O�`�F��ߑU��0Կ�z�q�I�ND��w�xq����PP4�d�n�]�<,���xI�:)I�ވt�|�o�7P��?H���cסMA�t%C*U&�m�����J�i�ONI���9�%�S�����y�H�֮v�IU����bEq'��<�"CKh�,��IM�<��NȆ�h1@p�8�D��t& tlg=<�X��ИKԡC��;���{p��!����Gڎ�������o������3��j+B�����۰�f3snbxU�|����3p���}�
ɓ%�I��n�N������M�&�8�ZP��eԸeذylKM��.B�"@���*'��M�
��=�CR��&�C��CY��5��M�n�
�.}� T�<!��s��(�G�f8�+���S�'e~���$�-j�yk4}s(�
��F�:���{�!ʫ+�D*6g����PTs1�5��l�uR�&O������d5�9�И�=rũɱg�)B���ir�{8#q�����3CX�{�f��M%�x`�'�BP� �K���lI�����9����_���9� SG�;���0O�<�z>�f� �]������D
�f+�����wEy�ǔ���-��'0��w���,�ʌ޿1�ډ�� ��d�	L��䧘],��|�'P����S)Q�;mTq�О�H��.�Y������Y�/�������� òu���j�b!P�4,�6c<ܩIs�6����x�ݹ1��ڎ��J�,� ��%���18t��E�&l�4<E����F�[�5^ٟmvf�2��˷p� � ���<��P靯���˸dG�>\w,�F������W�^E���Jx;��=���/&u�7u��r���A���|���ɼ�0��1���r4<�w����ƪ���YE����z��S}HYY �҈T��Z���/�:�E̰qI����:���h��;��OƗi��Y9t�w_ �|U����x�]�;�Q��<�?��<a�C�-����Ҟ���E�X�|Ę�{�rL����ƽ�����'��$v�I���l%!JU��G,F.�"�|P��i7<���G91�����-|Q��:�W����)`��2��ǔ������^�t�O+�X���xzY��1ҋ$�|ْ|�>3m��0����/��^��6	�(��V6A����z���������g�v0xY�X8
Z$X���t���Di�1�.�2�[ק�ݧlT��\���G;�s$ǋ�S	Q��2��H�	���Y΢e��}W=U�ߓĹ�	�oN4+��=Ĕ��}�Y��J�T궴%�3���x��t���]�27OQ�>�*�7�`0)ǽ���Jo:s���K��@��W�f�x��y�z90$�����ǿ�Ym�Z
e~�§�$�l$��\�
�lb�o-�l;w]>D�a&iMM��r�^�l^�	N���>.5�|H��o�.�� ѥ�}*����.������ɚ���-�o�]��&6�`�1��-��P]��k��.s�������P<�
���~��:O�6������.�<���?8�@W��@dg���n�F�{vl�b�d(�6l[�h}�8#�O@K��� e�'���$����-��M�(nv�b�"���R�[�~���gCSQ�Qsr��� QpL�S*H"�5�g�)����~����wlHO0�1�yZ��"F���@�'�o��9�]�o��Ij<�@?�Xyd�A�z�HF����C�����V�"�tч�ͬ���)s�n�g��6@9���}����1��	(�-] /�Nk
��߯n�?�!��8QL���\�dG��xx�z;��L{��aS$���|�2_֛޽��N_��/��5�o|=^7iz�8_1����f� w�#4��x39���z�)a�ڿ�$�t��wH��ƈ�7*�V�(�.Nn����Q���b[���ӿ�w"��.�vP�w���]���2� �v���\�V-*,e�=���]�s� ��8��;�#|�fߢ��t��;N[�C�ݐ�ܠ0?`�Ƌ0�wQ����"�M�<K~ޝ�}��"kn:�*-�'�����Z��5�����/���;�S��u�v\�my�!h���H�Ò?S��m��
1�����-%��v��>���0������q��֖0�Y�X.��f�{���N�%�@���"0n��_��$�V7�>��&����u3P�&�w9�I9�{�c\>�s��4O�·C��W��Fe�U!�V����Ȫ�av���GHN��T~�����g�����R��V��� ﯚN֝�v�7�</�=#�!$�[X���?�����ޘ�<`CJ��ú#�31Z�nD4�a���1�����*h�>^O��כ���K��^�V~�;�0�c 1`�w�Phi�%԰�V絹풦�����K��E�1�H�����W���nHJFUTk����0t}�Jn�EѸ�U��)�M4>�x@{` g4��%��xC����R��R��d!�t��c��d��["ᷱ�HK�޴ o�KM�uqK�� ������b��)�5��f{yK�b�K�g�j�����^��A�c��ȍ�C� H@���F���jѡ�VԀ��R���_����]�U�l��)��������dN�|���C�?�+G��9�W��61�jn�����V1�Z�G�ձ���hE	>C�ӫ�e2N���rw�o��s�RVQO���z�'w�]���Bk�{�?��=�Q=;����?��(Д7]n=H%�9ONϒ2��a�� �b� ��8Zi�p��^�v����#m�8�E.m)�Q�b2g��~S����>��evp�A_Z����r)Ó�?3z6�me���O��z��xn0|�*dE߇����0�r_��%�z<����#u!�~�;ۜ^�JF��X�"ҩ�v��ޣda��]��l����8t���F"�V�Zl�M;C&�9���{E���O��vjs����2L � ��7�v<��>��e��������9ݥ��+q&\�����V���7r�%�-�ѥ����ԉ��X�i���?Ü��.K�����J���ѯ\�Z4U���l�$P ֳ��O�O2�#�r9۬f�6��;>�xH=j�DR�)�h}MZ��C^�u�k�8��,l�����;Sߌ�����{�䟋EK�,�[	OSaGN_������TR�����S�@��6��Ow{��
��<�%c�<ޕ��|M;p#Ƥb���#�V� �,����+L�P嫯s��k��1a=,�JNcP>]��\'�.�A1J��u,���������/ˊ��q���o�.*/�co��[�Y�R��-�&�Vq�*h8�dcW����#Y��tX�ۂ�Jo�z��=�0�e
*&�S!�q�����$������k��4=|_��8T�c»����a䤒[W��Th=�}��;a�U$򡚘~N�HtRi�6m��ᬽ^c�z5g'?&f閑�OV���1�� 4mZ�+�2z%#B�BE���%��l���i��6�Iy�"�p!�W�b�J��Sܗ����ܶ6��݄f�i&��aõ��z_Hｰuzz'��k��6�9O�P�t��r%�Qd�|ƒAp����>�M���h��։B T�d�F���{|e�0f�$a��{�i)Rk��R�O�<wsYuC�IY�5P��34E�%X��#��9���^	�a
,s��b(�j%%�:��t���M�e���ݸ���qȕf�
�q�E�銘��~8���c#RcZ����QS1�YC�������W�8l҄gPxD����P2�6�+��voV)Wv�e��6a� �c���ܸ�b�]ƶ��U�þI,��>{{\ӟ�Ԯ¹��1)������oM�g��s�Jn�����^_mE���\L���D�G��s�wQz��8?:����`k��tu�8=!J�
��� b��3���KG��L	�8�z� �PK�t�lC>x�Ɛ�F^j������=�>d�z�B�S�0'�nm�2�+IU�a(�3�|��ͻ%֙�1qj�ƩW=Q�Zҋ%�A���:� p�]�;�v�}	�&��>���u��z��Ֆ{-���醦���Ax��U��_Ȅ\'�V��bu9�w	�Ab�u	�5�SzFT.�Ԅ~s5��l�O��o������,T%��$�Օķ���HA��;l�n����n�(hy3b��q��ﷻ�4���~G��2������ۑC��� �XR��	OC0�/nC$�I��^B��Bp���x1�JBe�So���Nqr 6��>!	O|�|�8����gN cy�<��D��J&�,B�D�iH9��3�%���G�61
'�e�T��
t[	S��D��=����8���N<f4���M�OFI5$mGx��{���R7�³k	�gϗ!W%��#��2C�0z�Zi�v�(y��z��/Wd%��@y��i°ȵ�ߔ��d�/:B0���e,$~�k��p�B�]����Q��Y�?����d����p h$���MSq�W�k�E�/`�;��TH쯂�N�����ǿ����S�Jp����+f=_����ݴ�Fzѝo�������:�)E��LN�&֌��{�n�1��M}����@��*1TƎ�,%���֍�]G?�|��1�p�z�9:��+J�b�Ӗ����G�Jv�f~�I����ټ$�v~ڿ,�"��mjs�����*_��N:��d�1�#?=|{�ڽu�9��e(��A�p����*�ۨ�����a�jv�Q;�.��7�B:�*h�mkO8�)�q��4�r�W����i8 @�	���\���{��yA��M˦�jDz�������1ʿq���=0�A�%%����BkU�����1�B@8z���@ԫQ?]MF��x���),x4�,+s��v�d}��G:�����@?�a/�~-W�OaW����s�����ϳ��$�:���o���h��9����g��&�Na����ho�� �ll�s���	�NO�p*mw�|Q|���`�� ���?z3+G5b�+6`W���y���
h>­N8>K�xJ�yQ`d��#<9�<��,��~��$/�f�b��Ts�P��^_�t�?��R�R�9�VB_�~?'G�(�s��X x��*�v�k�N�>$�[�pQ͚�D���ݪ�
�w�����܈	����품;��]h����N�2R��E^�������'�z�ffL�b��4�k��	�{}���G�rI���"O�lr��]�;��?8<;vߵ�
�Z{�og�˸G� Ѧ��V4���p�y�Ș��_���%����D��������{��2�5��{c=7��u��?9�F���J~8#�4TZ��z��)"x����_%!������aA�*��|"���
8"!��Jv�_�D��t��0���ņ�KК�1�֙z�A\�K�}�7�y��6����@Q�;T2�e��fM�	}7Y	U��UI���� *������BY��`,�L �ɇ&��i�}�e� ciu*!�\D�wԀP܀PT�6��1�'�5S!��x�,�gF"FiL���j<�|>��������N�q�-[^�&]&?R&�&R��N>ܐe܀�m�j~+�W��T�������+C�i3���;���>EقL�}K���p:��.
��K8g~���3�\=�����c��B}�$�5w3�9a���jOtc��p��P���
��s�p?�x�H��$t����k����TB�,��_2:��v�<נ�<��K�q3�見��2S�5H�����ʊzB�`M���v�F��z-�*����zl�u�=�HZM�Y�sc�����%�w]că�pb��D��s0D��`_�����{��W&X�y��n�
pdܑ�me���ٺ�R��Q󦉃��v�D2{xtq�u�L�I:�M�4�ޘ���A:�md=�s��s��Y�Y(nv*�<;��툚y�:T/U>ji����<�\��H>R`T3!��w�!�����d�Eb`dd��V���1f3����JJ������	���D6x����M�eVs''�b7�%��B]&铵$��6�ɓ���� :˺��V%=��)$8�5c��.:paϏ�6�K��:v�GgD��ms��;��|^����>õ^���6^����(�6�������=�������������j�g:�~ȊyDpkӃO�[�]�=X�r`�\��y["�m��zٞ�Y~�s�=�����-,AfTV��ʬx� ��V�5�����\�y~<�!$z)M$���w�hs?:J�h¶c��_LWߒk>�#���ri�<=/�:��OIM���T9O���׼�ZJa�NIH���o��r �}���xy�+�bEDDL�*ۣ�CC�cKɦB_�3�!��m�@6�n%��O*U��U^i)�e�������
�����w�.��HC�%�\�R��!�J]��XZjr*U��&���DK�k����^T'�ν��D.�k^�� �ũ����P�̭s����-��m'-�Eh��JE���B��㢊�G`��;gp������2H&0Pddd$O��\�`��g��[;=���a��]�X��B6f�ɕ�X9�,���B�e�R�]�.��������s�S}��h��#�C����འ�9�������n^^N�A��FT�k�?	���9|���Pbfw�p��4)x�����=��RP��(|Eظ�>%/kf����f,c��J�/����x�D�������l�#��2 ����=V����L�^����\�zNGG<�/�G<�xK9�ŏմ(�Ϣ��ClQ,���n���d.�`��ś�eai��Eް������s�3�=㯵b! �FU�Qn),@ӛ�\�sЍ�턌~�̑ܘ��SnC%���ŋ��j�v�:�`��$�U��-`hE`d<F}��X�y�hEc-hlą�8:9	ݼ��,=H%����z���|A�����!Q}�"A#$$��T{�l�a�jJj�F�`f�4i/$=��2�.P�Q!�e��E�z�No�Ҏ��Az@#Q��T��Ն��]`s+�8;-n�tum#$-^��m����>�ñ��.-�D�����	A}�HFs�!+�?P���K[�����򁶡���#s�1:X�����*���t�v��8[���!��3W����*^�k�V�h�:N�lw7u���oʎʞ5Y�ª;*��3E���- B���{�rmd���8����ZNl�t����;��Qҕ���d�B��$�b��!"� G���g�4~��2� �o�����\_qP_��[���^����HD0�U� P�1�>E����M�i�<�azT�����������Zo��:��;�!������e+	���[\��'[��R��ѱgg
���RRd�^�=�Dǔ۳S^��d��g̦�yV���������z�I*���8?F�)��c�Ϫ��� z�|߇���?�ump��8�r"!�p�ڊ&�Q!�wA]�{}�lm��:�6w���_Z�!��[>#��bʕ��c��Y��,.v[PQ �< | ����Bx��:_�Eb����S��B���l�jɭ���ҹE_����r3)�y�����]��N^�����ӈ��Ě�<%+��9���p>���������|��q��Mi,';щ������I^�'�^-'9"�	=JB�F�J#g(��d��Jr�mw�q~:�\��[�~u��Dӥ��y�0
R������Q�CsTf�^�(=+;��k^3�(�|5�S��,�^�Xx�};K�j�m]�mr���c5'�\m'A����P!����IE#��zv���=��[����$��������O.�^��Q$��J��^��	�_Z�>����U�)�(en̭��5��ڭE���4/9B���&X�˫�
qj9p���	xqo��At,���ˇ��:)=)��\:*�f�%9a��.֗<��rF��0��h_+J!;\��j!���1�t�����*!:A����!���h{z>���B���K쀱~2��c���wv���s���0^�%J��🜞^�_�u��U�hh���cH�~Wd���[I[Z�jؼ�������J��^��c��R~n\'$̯���!H�P��K]��C��'���Qo�ʁ�wfԬ�k����zRZ��9��_�?:"`�s���~�:GU �uѦ1�,_	H��j�,�����&��[��,�w:����aja��14�/��	�!���l_�^J��q�S�Ǐ���\E�#�F�-כT4ur��8�I��$W8�,�Ȟ��M��;ie��n&�6G��r��e/�/��:�t�T���Q5�5�P;4�sY��9��:��\��{|_s��~�5E��i�C%
�6vv�������R�T�MM��R\<<;p� Xؙ�ZYx�Ύ�ͨ��NB��n���&XBŝ��T*��ݢ�C��,U'��Tԅ�<�>��(t&����B�֢IJ8R4APY�� 6�����N���3�������"_M�-�v�1~�ų�B�{^5lҫUG���7}4�&e#�y�$�%�l�bC��A�I��6R�Oc�0Y1}�#�^�0��6����}>��|�   �YK+jaa!K�G9�i�����X��8O
?l������O����G=���|S����+�y�{��ḙ���T��O�[�kW�b7���<M������o��&��q tP����{4%`��s�W�"��Y��O�z�"�ݙB⿎γ]Z:c�o;�f]맏���!���޶���|�quh��z�[$x{�)��l�
ժ>]L�<��:x0����x����Ύ�[F_���,x�qp2�����Ip���W[~����[5�j�����J��YEv�a7���4%�R=n�F��s��/�#0�^9+[�ޔx����"TT[#�Wv��wGQ�E���K���k��ޱ�wV��.���c�z�~6b��΄体��Gk7��)(�Z!=���lͱU K.ujz:ddD������^�1�#<��-[E_LZN��'�D�n��:�_j	�!�Ǩ�w
����\-��ag����c��w�2��שIdX=��͐ֈ�N��x�T�q{[��u�V��mrPw�*Wj�6R���=F4m�7�q�W�G$�S�r#��Y�Ë��b�6������Ȃe�<>x���ł���'�j��e��ں�+�Z�0�͇H����36l�ʹP�K�����K�iψ�
L��'���ž��n+#�ϑ�%�_�t�3[�c]6~]�����|9�Z�	�+蹝�W�)�Ď��v��/����"���.���ໟ��L��p7IT����ʈ����%Ov��h9��x��p�K\�$8�É~(4��:aE�a�l\i����E���ՏO�;˫&��?1�� t��.f���@�vbUr�(��2)������k�1�c�������v>đj��J�y����]FfF��HxK���ܜ���t�:�P��w~�ӎ�T9F�n0�hUo�^N-I��i�x�b�D�`IO�3��) ^��Ak�x�d.�q5��nU�n�p�,'���H��{��Q���ߧ��1�I��Lnk'�\l,פ�0��q���7mH�|='��x~]�n��pt]A��\���3��m6����a2DvW�Y�dD��%���6����w���My_��6X؁�1����P�=����eh�O(	-�4�w"� p�|���.(��M�I9?r��"��EPG�@��I;�ů��� 87P���U�ڡ����=�c�6G�omaҾ^{]M��a��l+�¥�R-���[�$������nO;IC�7F�Z���]B����+���mwwww	��	�]�����ww�<@p��<�=|�����M�95̜3ջw����)������.�qs�I��\Ґ��w���"��h2�f��D�ӹ����=m.0�M��iæjQ�Y�G:)�q�FP�N3i{Y~S�6�z=�/�<�>_i��&2SA�{zu7�%�Z��]�05c��Wx������Q[˜�gFO.rp���r%lY���OG�ɏlg�{̗Ȱ�Q�}��I�0����|�+ɀ�_�̌�kt�"�Sh*�Bg�̣����2)*�F��L�  2�a�&�x���<�E��	����F
��z�Ϟ
O��<�J��9I�蚴l�@2��$�:���)4?tf�#s��rJ*nm�t_O�z�箿^]jhb�t��L�����~���u$�,�o���1���B������y�K��`u�������������s���jⲍ�����ݟ$eӅ*�Ë����-7|||1��6N��D���u��꺰�m=0��l��!�YOmS1�=��"�_r��p6��?�M�S37�������qހ��ɜKa)����Tbggګ2Ш�ÌW�X}�Abw��g"w�K���ۆ;d�E���o��x��e�M:%t��#�!����igm�����a��
�v���q�G��	r�|<[��lc�->I���C-55����8xF�+��?����Q#M��o��n�.v�5٣E}C8��U�T��8w�m��	2,:�[���}l~p�8z�P9��w(�yH;H`�DzTn���|�0����Bg��?Jb����e�˓X�y�`��85��_�p8l� w*��o�Ý�
'�}%]����I�f_L
� t�'��^J��s9��z�ږW����`�||�|�t�!�<�x���G�}z����Y����_?6'W��	�3z� ���%Y|� };,����Q��n�C߱k���Fc�*y����
ی�<7ڟ�����%>[�O�	��3�\�}�?o@�%$;��r3����>=�)[�}L��iZ�@�Sۆ"�#m�Rw�p���nIy����d�1w��
�t5�}�^��{�x������D@h�(f���;����%BNG���$P��h_�M��v~f�9j�y4�R���n�^�W����dK:|\�J��b)NZ��B�yM��v������2X��/�I,+_�i�n����E������6/��W�l�3����A[!��O)�v�h�s@��\a�>^�9/��(�e�H��u; ����|�5 Tq��E��B����
��J#��G
��z���ٟ�
��
�$O��F�-�*����MDjFw�Tm>�9���&>zƟH�0�w��$5��U�S%�C�� *���&��%�x�Vоb���T�X%W^�mj�k�cN����3W��2V�n�j�e����4�������(�Da�)��>�3�@A�s�^j�ұD��#�@���?���ٙ ���+��j.�L�/"��NcB���3���(b�:���.����Y-%̠rMmo�ꅂVߺ}ֆ�:�}��+��\5H:M�������=k�È���O�U�`��C��=� �Z�ky!��?	Ǩ?�[�����o>�;6겴�����:g�S���Q �� ��O����� ��ԸMm�/2����d�o�7�\��X�FI�.�b�Қ��5���&\�Cx������a��bC��L)��t�Z[I��|𶣕�\Ύ�P��iE>O]��!i�)��Ww��C��؉ �*F�h�?Z�]�ag'��m�V�#�3x�b��,E`歛<�(5���k@)�.�QqL�k_[��ɺ]�!>�)AV�X�k���r�HZEΎa$i|y�V�ى!�"Ob�V�>����mӣ
|�uj{A�Ϸ~"6���N-���m�c�G�����ⅹ9��B��r%z�D�����׏@y�K�(�;�5��Z����vϵ�`���r�AyU;~T!��`�ϑ\��!7���=�(Rk/T�%2�<lP}z�Ap�j��b�H����
��8��3��oM4�e̳�Ą�Uc��p�V������{�5����0�Nj��m9&.E�1��T��kyNk������'�z��#$�n��6�N����-�!F�󚠮iHV����e�,
���5un�y�L���cӝ����EJ�b����kZ<��w�"�˅��k�m]E�:�t�j���1ouF��A��r5MM8�?�$�LHX�5c"� ��M�&���X��Ҡ�|b��<��۟��fP�tx��S]���o���k}��Bh����'3�-������@+헝�e���M� �u%}������\���'c<���O.�x��!f���(�w�� u�}c��G27�IS��Uw��+��=t���A�,������	�W�����G�q�Ӌ�p�c�i0Q�O��]��о�T� ��md�\3���s����(�9m5��>IXd����Y���d�F����S.1o� $��|'�������w�Fi�H;�(��y�����%���������f���*��e&$���fވ�_�� x����Җ(��PNww��v]��s�\'777��,�zk) �	;��i�;�
��Ѡ�%N��J�}�v5�� �GRpxh���4���Y�H�]j����\vдXxt�h�Oe��Vs��q�?AN{k��iq�����+4nS��Y��ڶ�^��Rl�'�Dj
�8���?�X\I_>)����*}��K���}E�_;ֲݟ�N�|�u�w��v����i�Ae�n�,�_[�MY� ��*]���0����F�OvN�Xh͒"G�v#�z}�K����M}�x�:���:\�LޗF��g
��&�v��4ȣxq�p��s7���թ�����6��-�/^����o�d"H�}���0=/�ϊ�����[ ����o��?W$�/��O���qV�51�U��Cp[Gp�ى������A��=QB �غ��> B7����'�U�n=W����??�!�0)�ݸ5@�wY9!x�0l���1:H��l,�H��� �J�hn��~��������cn �O��M�4�3��5b��5�)2~,�	��`{�8��Jk"7��R:V;t�JW���B/�1?Km`Ѣ"�I���]��@R��g�S��۔����GE-�W�L4�z�%���z�����C$�Q��mthk�ed�[<�����4M:���H��7������(W�S������j��T%76J	:��"R��k3>}�e<u;�@C�eGG��3�;�ܖ��0����aa�Ez]A��ᛔܐ�r��%����TW�|
Re4�q���q@pl�e�͊Zs:ކ�u�!l� �N͎��FK�U�KIO�!���>�$R��gȺ�KL�tB��-+���^p-�&Rr��c����b
�[�X۶v?{���Ģ��,S��y�8)�u��	�v$�R�����<m�zs8QB��e�8�ę�p?hN���#!{�������&7%���zE,h�0�W��}�?�����.8��.�5h���3��C�C�ο�������z�ɩ"�k�f�2�!醾!=O���EШ�Q�Q���n?4�|�~գ����Y�r�C�~�]ÎF�{/�' ��.����-x��3���H1���}�_@��E���yqИ��+p�%��!ʏ�ի��}4��ݯ�W��>U ��)��v�o�z>c�U�W㑵��>]94�@��	�b�z���E���F��,��	�	�����I���T�8����`�?���/* �p�7B%�
D|t�&��In����ې��!r����{!!{�!x�4L�z��^�||��*�rz��E<ډ�7�Qz���.:
�<�ZZR"�����̃�O������ϳ�	絭nq֫?k՗>�c`<�M_K�^��'��vXwn_�d@�e筪��ϻ]���[m_ݞ���<�QH��9v�+�vW�����j�p�
@b߄|�A	��n�����f��2����@6����2)"ER�xe���;�j��s�|�Szs�C+��)��M���QZbk���(b&d�r��f�e|_������U4+x	�\X�W��X�"�.v�I��q٢����~�B./a�jp3M\���7�>�,4��teJ^�)��F~�7�5:)�4ut��D�#A��UU���F��!p�Yb����q-_�d^��
�	�p�T���sh?���`��tp1Po脚E���}�R6�SCL��1�J:Kt#O�~�[���E�ɠ�c5��2P����e������,�ාb߹�閭7sQ��!��Il�9b���A���*��GC$Ⲛ��� Bm���.H�P1RsZ0�b��o�J�@�)T{F��|��#��u�	ߣC��`�=�<��گ����6�򕶤D�^*�^y[|l��7>�͸���H���87�1�gd/����E�i�_6y����R�.��b���T�_Bp�4P�#Uf%$�r��aGbU�%!F�UoH�R����W�{K��8VX�VDL("Pn��ku�k�sǷ��Ya��m������BK|�Z���Y뱬(X���bnb�,�{Ǧ��ο�� �d�I)n°>�46�agt)��ށ�N�~�ƫr�Q/wJZ���}��W1�hѥ��EP�2kYfp�o�����^aQt�
<�U�	_�$%0�6�K��O|��Hγ��ư���n7X���I��Ƽ+�'	0�4~3��3K��j_�n2]�����e(��`"�s3�x��O��>�}���FU%�
¼�4�MT�e��䏇���q�9��*i���6����w�p�'3�Ψ1��N �P�g��lK}�F�����;  �K��	b��2���8D�c9��z�d<������?66v^{��U_�PbZ�v(^�*2e9#�h��Cgu=G�4:�x9�A�٧����ʋ�y�6�7Nz��B������q/
OF��>�B�%~�^��<�Y�=�|�~��E=9��r5.�@^Qu��{�Bmb�S{�/����O�&u��R�3s2�E���|k�sk\z޶g�Eav¤�����z[o��N�-�����Bo��y[f�N�L�/N�w�L�1}��;1l����r9�&u �Z������-�NN�C ��r�o�t�s��ح{�~`@�磫���:gKҿ�H�9۽=��i땧-��Ё��WZ?��j��9H�֬�������Y/M
�1>Np97a�^�IZ#�܂��)1��]߅\g<*�NF�i���ѥ���i���		��~2�D�)�|��O#�٥���g_p�!�{�?
xH�*mq���X	���ܯ��ٮ9$��f2vh<�B�x"o�&N�|����]H���Mτ"g�ھY��{t\�j��+݄���^۾{8lz�Ţ�����6���\ֈz��r`橰ߛ��a4���x3���w��f������|7��_x��Hm�Pj5LE�)3֣��bF��buQ���"��jI�t��a��jZ4$�_��L� �&��)@!��V���� jG���D��\W8�I�H�'O��J��P�k��Y��5&EJ5O}��XP>����4����GX�7�4�o3(=�<����&�ʽ��:�P�4/��`l�M�Ai����5��zϿB)�N�yWRKE�2��D���UA����!^�
��,�IL�U�L���AA�))>�:��O ͽj��������'EM��K��y\��z`i�]���jvB��I�H2���h)b���cU6�fI.:|���H�Qfǲ�ᗱ_P\`ɡ�q���J���%�#Ѻ��T�EZ38�����m���В�fu�4Y��;K��U�����<�A�V`5+�Z�Tq�g���-�0����|�3�%��sdddl�	�}��������2�H��� �/�DZ@�RH�_{j+84�vT'h�g�U�{�.��L���"|��O%b��R��x8$>�%��dUN���� _�y�4��i׉^����jk	K#���G���D����x�'����S�QP�G�zoTA>�S����W����Da�96>>�B�38c��J��P	
}��=9<
�P�E@΍�vƢ�w��	����D..[�T6��ZF��M�>Ԛ��30��/y���͸w����|�N�X�?��D���S�)���tݔT�t~�q�,P�_^M�d�q����p��Ɛ7�J�l�J�1�Fl΃���Q�Z�}sV��/��&���;�� ��V�C����A���֛LD�ԏZ^��`�v5�j�A��0��,���J=��>�I|^�]׿�49i #�yA��c�К�!���ԛ���mek29!��FWW��n-������d{�^C�
�M��d��d�L��C����]�[�3!@�������JPPP����D*����Y6�R�"�F-�O�p<�� ���ʽ�~������1��ߏ�@@A~��=�8��5��ɽH�w%�A���u�h�͝�s��8��Li+]گ��v\��Z:0���4t\9�e��y�;�!f"��n��Ҧ��M]co�΁�Qf�� IEe��^�%:���1���=v���P2�z���sR��,k�S���oi �7#�"5���yuS�����qk�h���l���b�2@Ĵ�/C=��͠�V�v%i�6�H�cه�Ͳ�� ��T|:I8��Ii�9�B^�ϲ W�����������#���1�s>����q�c���(�m�6��~����|�DlԈ��"��jw5f�ez/���;o�#K��ϊ�P��}<,''Ǆf��@�9���>8�6�儞�M�����9*﹗3�����������R��W��7�#���1���q`(�]��JB�_)�&�ƆtlJƒ�aLa�BC�\��$Zs#�s���9�ⵯ�3�Eޢq4Y�)�³6DTGe?`���p��ww+�����7Q�fЎ׻��1�9��%U%�1�ͰO����.$�Ќ�6n��~��37�9���t�w3�3�|���u�{��g���9�0����� ��i��>��i�D1DS�9n�!vc�:D|�gmm8���4�@�&Ad���dH��V���u�w�Avw�6���+	��*�Oϝv�ϞfV$�a�ӬT*;���w��3UD/0�Ư�
������-���a�������ׅ�i�O���g}B��G�DE�ϙ�t���u�)Ն���>���uKិ�	����ذ!�!���7�?M9��#����Ĭz��eк+���[��Zj�>f�\�9q>"�"|�`��UB��zOլ�#>�|�STDqh��������%��L
'ӛ�� /ݙQ`��������~?�*�Sd �]��KU�5�G���:�k�U�������?��!Z�a���Q��2/K�7����+(n��h!:�M��Ȱ�n����S:�_��Ϝ�'V������@����#�q��RQ���yО8�uC�NN�Di"O�K���O�:�q��ȟ��(����ơT���,����Դ�=]r�/(AHfFE<�����*3ȋ��t�<�la�;���XX��LL0x�������*���;!�}S�`v�@ Z v�U�q.����T?JL�]5|�d��c0,��PF��<#���� vX��w�\���=_�ؾ��ܒ5�ǳ;���v����"4��9@�	Qީ]��mJ_w��%�o�)�v���Dk� �DUB�	W����.ZY�0.������Ed����~ ����5Ʋ�e+�/V*�҅�>��2��Χ��v"u����8:x\����(@|u�����X��C:q����J;E�Ó�˱�]H��H�/��U�Ս<o�D���Y�t����t+��)Z{{;�W�do����ӞI2���7 ��כ���SnaM+h�wa{a��d+x`M�>M/��=`��|)�ʯ�1�%K����d�����g�b��ז
����]U�{PZ>?0-c|@.�M�%a\zVo���x�v��#��� �<�=�'�|�xUv����%�t)�[�Xֳ�~�'�I(����.h�64V+�XN�b̋zˈ�)���@!`��ŗA�x�:����`�;����贪���=�{���;vΒ�Z4�e���Lpp0drrr��<�N�{P ̎��zS�������Vq���PԿ�ݨ9B|���k��wg��3�TN�
z�-� ��7M[�+�����]��5f=60w�`�\6�B���K��y���	����w)%mIky���<j_ O��i�d�E��qU��@f��/��c��)����J����^$
���s��Zc����pq��Q��� �[�N�-|m
��x�$����<<vD_wE�nU�66��Ӕ($B��� #[)�뵬�VFCc��hZ��\��I�yV��>���b�Bs�ej����<9�P{|WP���B�͓�ǉq��9p9�5������\@O4��^�(�� <g k8�˧`�i���j'����)o?��(RM��f��$:����㛗��p�C�W]Ԯxk�G�n�����T���Zt�l���>�#]V_�hFae``>����kyz�{��v/���[��U��5���#�Ѣ�ȡwvv|�?](�����Ϳ���~gboo�ߛ�h���+_V^.�.b�����΋Ȅ)�0��|��X�~�p<-�Q���#پ�d�xr}E{P���H�ɱWH�6��Wi����'�$�Z�({#�/����!1�F���_���A�5��'>�!Htc'S�o�J8���H�)/���!�Tɸ	I���:�
z��ja��4����=};��aז�^~��V�ᗃ꒎�u�}���(L����Is4�D�&3\��%�����zZ���ӟ?�^�[���u��8�Pz�y<>2[4�8'd���c��`�a>]x{{{e��WG��!�9sF�}n�}ؕ1�Rh���BUW:"��X��A��d=�3k�� tLZ�${�8<�������F�E�)XhB&�'3�q��H�a�[�
M�k|y���54����z�������>�yv( %�؝cys���z�����C�����0N��sT��:���'��Y��*��GrYQ�_1��'Y���-h�R�����`���.j,$����I�U�lD/���M�!���L�'F��o��2B�u���T���j����5D�(ihH
HWNc��,�@�i=�tH�r'v�!�s�5�%�Y�f3Д���f��/>yj�&�8}���}��f���A�Ű�bئ蒨���K�sy�pB�3:���?�c�9]B�S ɝW6Dյ�:�G8��U�k��B#��>k`D������r't3x���c�������9��.�G~�Z͙����ɟ��^0��l��?B7\����/Y����s/�Ϋ���yd����:�.��10��Zn��ۓ8���F�3���|Dݟʍ�����S�u���p`;إzީV������	�Ԝ��w*�t��:*M�ƀ0�>��#�+��-@n�ED)�郵��v�9gU=ږD]y	�]Hl����g2�N��N,�QB���E��;�]��=���dȃ�,񙲑���Rj.PpF��5cr_N�����r|�����׶	�b�ֿ��٧��!/�^�Y��n���â>T�`pbbb�n>Eh����ˡ��(�O	�i�='�?Q`��D�2��ǑE��ڧT'7Pҫ&�h@�/0�PZk�<)�ӎ#7Ð��s�b�(���&"���� �6��'3�~_���U�,��h�f�!����8o��`!墁Y��H���X�Gd3o�eA�Tpq\���f=�j"�j	���4B�����{8nr1�4�.�����#��V<��s�9]����O_w�v�](�S�[���\����P�x��f��w�VW ���� Vw��}�^a����DJRF�n�*�0Bz'p���s��}�{#���)W���S���>p(�����;�k�%�<���q�œ�kz�!�^�8j��6L��*�����Q�W힮��<�R忷�K�Ka���^>����G4��lAϝ��FC�S�� MDFA�sh ��?�ぁc�l�����]g�$�����'���M���\�:� �1��������$��O/º׺�[H�]U��q�5�W��V�؋�,�tO9ִ�c28��m~2Q�"hHl���D��r��	/��Ps�[6E�c�����f�~��@�5i�u~{�7;���s�o�w�A���v�Ǎ��3n���Y7�>��MM�fQbCet���K�1EB ;��([}ٞQ��<��턉���)))��J�0�<۽��3�I~~yYs�.2��*f��_m);t�etl;D뉮�U�r�^�ȺsV׃�I�M{�`��0�k�t��ž7�'@�߯�ds�y�T$FR��*J¿�L$����E��%�B�N�1��_��?���=9������R�ԑ|�b������ѐ�D5��M��nGjU������������u��T1[B�eڟz�LDQ�ז��z��]ҡ�1�Ϋ�x�tʞ��_�����ڙ��]�v	�V�P|)N�H��<��p��#q|�d��2����t�gl}f*�j��X��������gE�%��Feuu�a�0q��W �aX��Qs�>c�f��p��:(7��-�w��59����JIO�a�"��^B����y55�>| ����S�?�ճ�V��Ċ�z�\��/�b�T?!�rN^E�H�Տ�a:I� �i�40�@~�Xŕ�d���Q�hs$�vb��Řl�e����)�w�y�Vg����K+�HZZ�K��j���3�X�SѨ���1��j<�(�u��2��� `������<����4�#FM��)h�T�x�g<�����!���)�F��!��z��Ly��QU%+M���,py�o��,3mS8��I��JU�?=�4	�8��"zLZB��W�:x�������q����^����i������)G����g�I�55!A�5�8�%S�+*T4���p�u
��-�UPPf�b��E�:<��(��jf�$�/���a��&�Kq3�����^��Z���6������� �u3�7���"����$lmTg{�OG���e��Z�y2�y�_��Q�q�qwx��$JB����n�+8�xՍb)�}�gT�F��k�>:w����Z���������w��ON�>�!�k����%�A4�=�����Ynn���~"df����(�#���؍Fa$o&V�3�	F�َ[��9���!:
��yo��y��0���|g�3���u�*�N�a��>Ƽ9/k����sS������3�ǁ�F���Q<h�.�=�nOX����y���;�'�{�	�u�]D�K�\$
�e�K��Z�*�z��j7! 5l�n2��ď��^;>�i���21_� �j�^ ��VS:7A^��r�3�7%�?}[�F8\Yʺ�TK��;f����a���%��5X�C)��{��_p���)�HG`��S�ۖ3�sE��[�䷴I��������Xtn���"�s<�҆��(��|=Q�!X�ń��q�l�����5C��tn�b,ŞE�=:�]��:2e�Qlh$�'?~^�-O�CeK}E9l�z2�~<�j�z#�jopF4fcbddd�^�J�_@>>���=*?Ñ��tzG�ab`�:;C�
$�2Q��4B??�o3��`�����4��E/8Y;ڠx~Qp�~{�#][�s��-v �Ƙ0F&��6;&k�b`L# �||�F���U�t#Q����ǧw��:{�y���-KjXtʂm�liv|�c�P��&��Ev��	��&N�ay�o8��*n`��.��#5ޠHxpn�I{���`L�Cx�����8��@�/v�Ah<��i
F��\�|,`��S~:l�T��%Pr�*&�:P�2����ôQ���j����[R�	$%���$͓+Nc\I_n��me���xC"��w��)����,���h�Ca����QW���8bU0jfY?�!:D��������=������9E:ં�H=5U�R3�>�����`�ʼ�N=�dO(ñ	��q �RkW9.�4]������r�����f�����e@W՚հ�i&�nEݣ����{��ڌ�2읙��������^v�)�9��n��y�h��Q_�-(��fT�5�Iho#0��x�'�n�إʦD��L�:�Xr��GHt��c�U����Z>V�~�ན�<�]E�K�r��pi����
e$�4đ^��K���js���>*�Wڕ�B���w�
��I8o��)0*���1�t�eX��2�$���/4�t)�K�_q߃5sJ>���.���������jXW�?�>�D�ؠ3t�(�"��uC,!r맰��
���UH��,F�g��\�R �Bk?}�ܓ����|�N�������_��T��o�5ۢ�(5�'"�t��U�[if�^B-|O��~�?�ǊzW��AtX�j��:��:��-������8��׵" j�(���Y?��鯇�,H�g��� -�����˞�j��Q�^M������P9����:��3��vG��
��*��r�ݦ�z�D��;V�.�ipl�R�zD��΅�7�tD�w!GH,p�eT��/v@}ϸ�O�nk�L�&��?�k�S?7�}<Ԩ�Y�XdN����l��-:�����<̾�"��G��%t�;r�̇�fp�V�oK*�b�;.�7��Rih�Ǧy*����_j-�U�@,��H5K4h�3&�!V����P�ˀ��^��"C�Jo6xć����y��Ҿ�~2mr��s�^��r?0OR�-�ܤ��;��9b���Ft�$�\��F��@L���J�M�JC?A��q/�7�7���6�ժ˥j�ء������*����M���	��_9-�P���-/j��v��Ư�����Z���<s�kD(�@��p�:}�5�sE5���\"z�V�B��éu~�Y1dTIj���Nv�v}�f�</�nO'8H��.�g�}�S�6_�L�Q�I���c��O��;��=�:k��Hd���x�yu7��;LKe���@�TӍ�۲2�`�4AZ����~�,�;=��Ǹ�����%�	�x:BZ[�.�Yp�Y�#c'[�L�/AJ��H�g!%{�޴���x���	�ZF��������ŧ�2~	|ݗ;�Wq���'����&���)�=��&숃˺���r�������kד�����N�;�<�]&]��kؕ�������j0Mf�Ө����o�+��_7"�6ɪ��>PxN)����z���=�W�r��<�:�:�N,-��l�V����.a����ŇCR֭]�Z�v+�2P<�SGYƕT�����d	�#�;<s��nu��/��(i,TA��P_	��y�jV�`9(�9w�|nC��7�깂:<�y�����F_zot����(�s�a�4iJ9�{�C���fe����G���;��W �=s��o��pD��{q7��oGz��>\Xv�zY���i6#��6�}M��7C=�X�z�i�}	�L��C�,�.R�@��I�"~Ґٰ�s��mU����:zh�������Y�Ы�Ԟa��fD��$��r����}�*�~SQ�Ϊ#� ����9�(w��GU�F�L���9��'N�f������߽�����[�ڝ5�CPX;`N5�b�㢻u�ek� �*��;��%�����j+��z�k  �����/M�a6���U84.��g��/�{=�	|�6yF#w��2z\�ş~�T��R'��I���Pz"�AH$�1�H��/�8,ںF( �����E�O�)�^�6�U�	�;��k(_�M�3$J|e���d�[NVd�-|]k����u5Q����s�)���P��;uD��Uj��5��v?���n����ا��[�RS�7|A	��1k{Cd�ޓD���s*4L|خ��q�؍2�cC�V�y:��6��+����k>�b�G��)�hh$(��WC/�����Y{�,���)ښ�q��t@Xkf:�i�P]{��o{�*:�|@�?��>��:h�*�v��l�h����cGZ��տ 3�'�,���F�Q�ۼ�����x^�p���nE�8���c�`m���Y������X��C{�ř����[�&��T�����틳X#�O"��%3��+*X�㵩�ڿoۏ~����5b�`D�U�������<:���[�x�^�{R��.�����ѹ; p�o��5�����WO�����Yv1f�_��,Hx���V�f��������x�tL���2-lX>x�W\�^�M$\1���>&��J�L_l��&�f�'1$������=�P��0��~)]a$.c}(����ȻmV.o������v��#J�!����:��M�o�o���||	f5n�B7%����i��}Y������iv�MD�7�O�V,�Q�4��mڢ���@6��wֈ$D��&Sjm���1������`9�S��l���1�g�'���4�$� ���wK�y[C�~�o�`[دܱ�~�?��D��y���j*vԜ�e�t��8'��s���J5~��޲=v\���~uI�K֊�O]@����u���G��$;�x���_�!Z{B|�������TPK�$����΃�y��d�i�:��R�O�xlwzL��S���~b8��]5���2P5��b|���Y��lX�ST_K>A�Ɂ�+�
]��f�
��FdK`u��|
f��hg�B����l���E^_7�[�\��xz�H���:���^j4��k���s�g~f`N��Z�^���´��r�G��JU뾢��D:S��;{�4�]�B� �3���p�[Y��&�j۔Q����O�VyT�yt�e�x�x�jl�3F��{������ߥ�s5ǟs��	���P{�ޢE�c��9Mf��z����f���/�[+p��A��Szaw?��A�pa���n�ƶ>���i�V\����o'�k�E�W�&��e����)N(�d�Q�rL�Gk_5s�iI�=}�載`�`�E,�N�%��]tw��矶��Z��_&8���<g��[^@5�I���O~�t�6O��찶�\��=}���7����uq��o߷t�B5�z% 8?_Rk�}��)�c�ZG�1�����`=̇G�\�=6-����"�?���[��ݗ�h'�/�M�_B�h�N_�����A���Uu�T����"
y[Ջv�iI�w�b��g�堙���g>Oo��kM>ʇ(t�����t9^�"�k�52�o�y��?`
�?�q��K�)��S������.&<��0]�KB��L�Q�ve�Y�����ԸC(5�g��Y-fTpN�@79������xg؉��%V������6�=���h)XǢ�=��*P�}�ir}�$b� ��e�\�3a�ץoG�/�R���/�'=����9��ɓ1l��N�X���7SO]��j�p�6�j%����2�T��W�?��G����I������bF�nzH�';�!Lh�i��:m{�D��M�,my=!*y��x"�v�/�:T���,�;����4���YҞ���p6�mo���o�z��[+��˱�&n^����M;���/$0��B�b�C'[}�.��Q�2���πS��j#oB8���N��~�S�p��xǒ"K�p�M����XjD�����6̑[{�Q,����M�����<3�\���@|����������N��*\�(������R��gC(�J�3�d9�T�~�U2�l��/D�?�5w �GS��{x���69��۲Vdol��d�qS��P��RCX����HW�o8�7�=*	����W�>���b$*wpr�}_u���QE2-�Y�z*f���8V�Q�&�f?���OǗ���d��4�Dsz�%Ζ}�Af�_/�#�S����R=���+���F&��1fx�YДe��tF�FĂ�/����:�ܤ�@=υh�FF��=μ��6O�r��}�Z<D8�S���5'Th�3-��	�tǾ@�d����LpWD��ՙ	��)k�H1�	m{��cWr�u_{���N<��+6�l��xw�[g%Y�k.�VR��V��&|�<d�Ώ�U������D-*1�<�,#�7�t4�y0�a���ʲN|u�lI5��lL��~����ͭO]	���S��>��V��=E��m�Z��}68Ǭ6L�}�����a-_$F�3��W�Z�g� ����+-�T�$R&xH~_�$�@h�!iQ�e�Z6v3GJ'좊���WҢ��m���{����-ܠ����{�*��Yˮ�:�)����Ӊ�?��K���芡��ۭ�,����� zy.�@� ��Gs�+C�b����[�hf�x=qZ��^]�'�/�$����}Z�_b=
�I�ژ,}{>`���TT�cnКɃʿ�|n������L�R'�P{��o�]_+Z�AQ��7�ny��s���t�Ã;���!�wwwww����݃�&�������'�+����a�T�޽W����>5��b7���Z?g�켯>m}�$;l��G��qo�O4;�E#>��r[>��w_�h��b"�Q�C [��[ٻQ�D��⯖W%��u�n�h��	�O���G���D�Y��R{ �,~p��۲���z�Ğ�W,]��=w}����{�f�W�]Ix��6���U[��5���gN�!6=���D���\��� ��O�I�@ű6y #��n������60P>�wt�F	�!�j裂(�P��;�D���ި�������\Kџn��,��u.]�q�f=���=7�fQ8@D��A#������t�}rq�U"�	��1�/��a7����l'�3�_�ZGn{y؟?H�}o���u���@�/B$<�r�m$��½���Ih%ڳq����%�ɢK�43�m�y ��+����m�v�/��X�Kc LS�=���hIG>Ǹ �j���>�Vs�����-[�SJ}4f���w��ݬ�00�&����ȑcH8}���B���&M�����&D�9q� �~�Ȣo*j�Y��df׷�K������zv�:��]יh��!�z%���)��v������p4��<.��YD@E�(}j��y�ג3��s� ��d0]�q��BF�tq�XSe�s���1a��J~c�'�]l}�=�jh�(�n��j� ��c ����$���,Z> r�Y����m�?�l��3���$ad�;�aQ�w *�e�>��Z�� ��~R���1|dr�}�)onx�?��^��Ȼ�T}߽��+]���'Տ۱�b��s����!���m��(���pZ�u�e�H�9�W[�F�P�������JB���N�3����7"�I��6Cn4y��n�G�8�|�y��|q�a�.�y˸'^��Ԏ��{��о�VB�M�hb�`��}2�6SU�u�1 l4��h��%�{�>���2m�Hc�l��F����F9+���̲����d 	~�̫�3�"ȝ08/�Z	���ʱ��W�OZ!.W������W�Y��I�f���H���@A��T��#iz�k�t$�����eVPh�y��\ �%l��h$����?V����	�j�B%4���z>�U2�M��9��XI��i��m\�x�:����Ā0��m�hv����⺦��O� �]&��~=Y��f7��X,�:s(��&�i���؜��#��:��"�*ǫ�OK�>�O�͸����ZI���>J�݂@5�x�6��J�^J�\�K"�1�e�M�
c0_�j3�^����V_�D�	S�7J�1R��ń�]&D�q��ڥ��jrw,��t��|�r�������sPҎ,(�u&�	�c�DM�j{Q`���wt��a]i����j��[Eؕ��+QVÎ�Lr$U�~Qm$΁�V��U %"3#��o��Q$.�Ly��bƠ$@��2��l(!��a���;�c;fN���}��'��LN�ciwÁ�������@G��~�jO�7ƚʬ��P�>.�_�r�j؈yz5,�͟Vw����$�{�T����Yߖ���,#"�l��m��2��o!.�ӌ��G��,rOW�2+�P���jԦ#�V:��j�zЮ�R��}��&�(k���k���\�s����5��'_i��Y7�mI�R\/9�F��>V���>�P̿����x5��	0�	(�{w�$	��Go=��*O�y��>j$	`9�"M��̼p��D�ˋ Q�Or��QR&���3�â~�p�d�V� 0:�Bo�[�h
>4{$@'�F����|:�>:V8K��{n�׆:g>qz�By`�>�^a٧+�q]����[�G�GM�IR}��G]8Tl�����ߤh(�Q���U�"a�1�F���PB�p�e:+q�j؅J�����Ћ++G�
Nf�Y�5*�3<&��p_tɍ���U�*��mMvS��k�>��I��u}p�
n�Vt���Aa���]&Lц�GC�:%d�Y��;��˷�������{w�z�
��O\ywJ�o��3f�������#���#���pj�Kt>��f��\�P�X�L���zҥj���YY��1�,��L�4f�cG�͞��!�7#�m���& �`?)�!ڜ�1?v[�,�Y�Z�
�<�ƴ�y�:t�7��/8k���M���p���**(��CF/�q}���O�)ID�M/���Ǜs��A�&���Jo#$�]��($	��ݻY9��$���n դ�IE�sC�O��q��q糶�49������� ���9�?0���x���������z�N� C�Y�p�����I��~{wYY���r̰qд�-�K���F�ۥ����ok�߸�n���ͬE��k� b܇�%!��OIR�ifb�]� M��F��c�
�T�fs�$@�iXM��7T<>Hy�2�d"B�.T�~���;�:[:�������3��$���H�Vpp�]H���=%wOFR 0ٰ�
�u�yv7��j�#J��Ng��I�st�륈De��ԝ�L��X$5���������� 9 \�X�
�Y��0���})�++D��/l��֪&̡L�Ύ����7� �cD	;m�ޖ	w]��)��%׍b׹ݣׇk��
�\��e�� �@�Rw#33Jq��Y6vv��Y.;Εxq
J�Z@A�p>�|��g��"C
���#@�<<��-2@�k��y��{�NdEx������=2[��>�"���U���\�;g=��^9p�.Vn^v|��U�*��v̅��SU�)E�$.j��g,Dl_�|������(Oxb?fL/�s.�����jI��=�����S����9v��1�~C I��uWǷ�g�ӎxZ�����fe %�����`Aj�s@��8���&��#�ƪ�pnC���tQۀ@b@�'hȓz����_�Rc�����\��6��~�C��6�7jY����\�0Km��^���o�FG�'@`��~E>2�U������n����?�;�f%,l���OU����_����T��~2����'�AG���Kf+ʣ�ҋ܆�cS�����I��%����j�f���������1]4d�N��+q
����&n0�ҙϹ|sӃ�̹�tQ��V��W��>6\���zCy7?2�rn V��?B�ў���aь��E&͗q��]ӫ:�@��5?	�I�L���>r���\se����q����@E(�`Xf�J" yQ��j $u�}_�t����QϏ���ŝ*}X�H��e������&z�eii|2ev+`zj�ב6���j�+�έ��vB�iw�&��s�ᣀ�H����'�q��Y�A��}�YXu�Q�v�;A�x�Y�����1�f�+\ ���	;,ܞ#��+�˶�}����6�
1�t��Z����M%�d�ڷ1:���2�2�X�W�#k �UO�rjk�*.�fJO�
Ñ7W"� ]�0�k-�= P�?� � �O�=��O���cwY��6��̗���R��V�Kx�h�[=5�Ѽ ���>�d_�+�Y����Mӄ~sC����<�:MیnÅ�$��';U�����y#6$]t�8��4kP�R-j��g����PWCS�����;�����l�<V��vsJ���b�G�)��h
?����MU�)r��P~92(7��xbOԓ�7���(0��2H�|$�Җ�i~�����^!e����	566����O�~fH)P��O������V��6�����@�f����Q]�ME�ܑ��η��L�A�<�Rp�Rm�Q�@�
LQW=I�T��|��y�n�����yk)v�i.&�s 󱷋���:�������tA3��8�>!*�Ĩf��p[�J��N�Ξ�͞6���t�3e��#ƚ�T�I��m�ًf�v~��C���w=���Ҧ��ug�C-)݄Hv?SN:_�-�s�Ud����~O��ܞPp��z]�(v��Ŗ��ǳ�s*��<��5����4iVm�5���'�����C@t�JA�Ƿ�-����NK�7׭���Y���eS,�@����}��$3@�p�_Y�>����5�����5ɢ)L��\�d��3ڣ��� ��ᷴ;���0 r���,te�N�8�}?���5�0�5�2��} �=J��y=�y�b��vM놻ǡ*e��#����M���J�40�	�9�4�žzt�A(��!���={t'�qfw��{��M�
�-��_m#D<?�1��MpTE��44�~�`�R^p��I�w�\dB~ȝ=�Wý^���c���!��+�VQ&���bv�1�����#b�,^����t?�ǆ�&�a���K�WE&&h�l5����U  ���q 9U_�M�`
�ؚӑ��'�]L�'aU��f��\�����*�'�2\`^`$�w��>:E4u:��-�L$�F�--S�6���z��~���!�A��=����)xʴn�ɕz�����0P��I��~��˥\�n�K�4���`� ��k��e"z���{���'��͆zW�A�]�N��U%�O�2�Z�Q��(b8���In17{�1�G���_ T�yB�8o�L��s�g�!m�B�����Hq�E�T�_Ru��t{!o^����ե�G)Ä����BA]+A�Ct�M2pE#FX����(~�˴���s�bQ�-���׀� �
�����?280[;�c�G������
�h(��p��D�o��2���U��T���T��)�e�P��\iݹ�S�`����QN�"�Ӕ� y�ڇq��җ��ZDT� �'���őۏ'��� �'�L��^XȄ��cFQJ���5s����R=����	-��~@]56��.���bd&��(fE���Y�@��F�@ ���UƯ�#�.j@��
&4���w�߽c;��˓��'-c�w�a`BDb,:a�?�3���y�W������+�*�'EJA�6dEQVW�a�Y�(�aN��j��*�~d2�t�h�R*ּFV�W~q~�HOvx�I7��'v��i�0I��`�U��A��7ɿKY ��q��~'2E ���;�EM{3��������&{�.sƮ�e(��@xT��@�C������;��4���SI%WP���F]zZ�5L�_k+z��N%~�3A��[�8�{M܂�x�k �¯2RpJ���X}���XW�d���e|+�W�����_w�I���/�=B����˩�C�\�*���ږ���by3�œz 1l�@�4�@%2Z�a{�|�gU�}]�ݷ��$D�2DD�;,�D&E%�^m��wD:��u��m�����&U� �'K7�����23�z}5�h�(���^)]��[��'`����{����m����9a�j�՞�����/���/��u��-ϖ�lQ`��|���8��9�x��BL�P�4�.�x� ކQF�JN�5�U�<%죙U����]�"�� iN��C�5�n�u,ځ����.eD�˩���y�F[����OV���TM˄ԎO��]�7{k��T������Z��I�4{�!]�7�k[s�M��0Nd��/|>�k�G��1Fs�Q{�&\	'�
����T���&�_����:y���:�9���n[��t���5J��a��dS�XǼzA��{��Q���!!_��?����U/�����!���ҵ�U��Ϯ�LmQ�ĝ港�/�T�ZoX3�h���M�
�(��V5g*�iw+��Ř$G����P��F���`t>�`��;����A�奄�����t�x5</Κ��KX�z���F;|9+���*���f��	k�e��W�2�Y�ʺ>�Q��x��.+ף�)
D���Sz�����fP]�=O���ּ�;��1-�;^/t����W��<�w�=`"J�4��r������!BMA��B���������J�$w�	�?�iW|��a�kj�x�j�EX����9>�������7�i^G3��i]�0Epeg�q��V���p���փ��%/�:[eg�<��;�o�7�1�E����_e1n/��5S�V���*1���ԛJϹSB_<喚2�S�"��>�!؂8�9U:Ci(~DEZ��V���k����W�,q�R$��u����62t?����Y,�����]ɐ�e��u1UW0�m4�QR��������k満�/R���	�}H�H�������߀�i��Q�d�0��F�"
�L��a'b1 ߸�|�C�I76Ҳ��N\\շh 0����qft��O�~�VOar��Qj((xtt�Y�=���H�Ï(���0Y�D##�9?:��!�w��������kr�Y��
�������HD����u���p������~XcM��ˆ�]Ƣ��5��k����v"��5uT{��Q��_4č��:CŁ�I^\3��b�UA\�W���0f_M>y�_�c���?�~�byRc���Z���_�m0 ��c�hR�~f-w_[���m�βC ���f����w��z����Dx�4��9�¾j�,�h���a��`���pH(��"8i��A"ZW�*��&7��|��Q�D����L�23o�D��M��D=�xFˎ`��N��Hw��8��<�B*�olɔ�PT�l��Zs/�0�-�-�}�+6�-17�ˁ� O5	H1��B޸�!Vm�+�]B_Íᱟ[����o�Y�5��o<@�X��}@s?r�ˢZ[3L�#y�hzV6��.�`�c�NY�#)Vp?y�豂΍L�K��8%:��S�\H�l^IЖ�(��Iu�6�f����5�`d�JY=��P?-��Y�ym\��R���+\�O|����x�x���"����p������o3la"P�����/TQƽHIΣd�W�ح�Ș�1U���Cd�e��� ���`�.x�B�U_�b�9��Z{����y��z�z�.�d����Y��@�?G
���u|�VO�CUGЦ$�*Y���}{m�����[�ǂ�;�5$Hm��ڢ d�}�>D1�,`6���3� ��(? ,�h�hvˢ���F�e]�aH�\�������|�,���
maaS��<y�IU.��������0v5_���ݧ�d	q�9v$R|drqӒ�x:A�� Y���1��(u�R���.S�:��Ҿ���4W�Y���Cl�EVF
�U��^�,;�a�����"e���~r�D�X�E�0x��1Fb��xvA�	�֭�&�R�Cʫ�I��ԏ��C���h(J�<4?�O���,�t�90	�,�3n�SVY	�f�����v� ��͏+)��DB��:�0x�s����хQ1t+�V�YVl.�4fO������RQe/�w@��2��@�ؠg���s�s��|Q��y�PɊ�w^9:�ve��´�2z��2����y�߁���9l�0�K؞��
˜�,���ۈRW6���:R!Rd�qqj��IX1x�ߧL��PN8#o��AV3����4#+}��`�iW������ks��z��L�f��PR�A�6���a��zl�1iۡ�[9NଔQ�?�
6�0cL���y+��I�jd<=xTgt�	�XS)�����nI�Ľͻ���(�P�X��DF&�?���b&A\=���S����}��4��s6ZA@Cq�����S��~�ȧ����}�y匑�"K���䁫�P�Y+�%y��gsU�,y��'W���	^���+]�A�s+�(;@h[��5�]��-����[.����
����t5��a(CL�^'��	kL-�u��$h��#��j��g���:{�p��h��?�ׅ��P����kIL#M1�Ч���g��[MG�f�:���3�����]���6�<��E2
v�R@�;�N�4��~�WM9��PK�qG$�u���0@�`3Y.%7����zt�yd���-'n����4bO��A�Gԝ���*pG]�tD�a
P8:�@����ɤ�mg��@)U��	�^�ՉJ.җb3ԟp���5����[q�6G.�6�&����ܔ���Mn��������M�dV�y/�E�b�/t9�$W��Fz� �+�=�I��v����H/����94�TC�}���i������{��G���6�{`�|��W�	헠����!/"i�c�>�*Z*�w�%Vk�
q���d�L��{p�n��`Q�C���4��dɠ�Q#�{�s]0YA�7�)!na���«>r��bG�KX�.E�~�1�+ �O����͟j��=&�j�9W��D�|7��Ф(�����s/t�
NA�9�S���)��>�[�lu��o���ڍ�bo�wV�?o�/�{�U�����z�.��>̮{���5E��n���"7Ҧ��r�#�#Kj���韖���P��u�˥�H�v/_���uh����m���t�`hP)�#�]4�z����{<�����8���V�}�����p��4��c)5���HfQ+r(!�J��</��O��?��_��;��
퐌��w��J����i��.��H�X.z�<���U͆���y�����6	��m�K��.��NGc�%=��u������ �t�%7A��ZÍ{6�Q
z6N�`����@�J �E}�L���jӛ���,�㬛if�I�T��Z]tb���v���×��ڶM��9����=��{2$�����
)��|L	�_x�8�ѷ[9k���Ev�M2�h
��-�5����Z��KpyE���t��C�c]��}��� �A��/�>\�����C*S�ʯ����)�;p�~m�A8u桝�6£��W�Ȳ������T�t);z�,+��O���������SC���iנ��JE�l�Q��9޶8��{�wͯ~]tf[�e���f	1�^�)�z��'�Vm�
=@^��g�P��6���^��c�:v���kt�~$7�(yE!�$�4& ������K��(����ӳ1wo�C�}�j�'����!F��6s'/���FًJ����_��	��#���7�E| p���kpr�ә�!<��I�������8��R�v�b/��N��p��	g��9ݔ��BW��B�-��jQUɡ^K���ij��#��ֳ�掠�i�P'��?MmE�ɬz.H���{
&M!V�Ԁ�
�ޤJ1�Ox��y]윪��o܃*�q~hu���G���h�_��s2��I(G�~]p���l95g�ѷ~�f�Ao���d�}�����t��Ty�d=i'��
D�����~�Ot���m�5�3C�0~�Ӡ	����E_��q���������J(@X���C��Q��������э�RL�{�pR�?�m����z�	F�l�<g��Y�:b��z�,��z��ϟIٻ����W�l
RfC'N��n��l�O�|q=���9�'�_(���x�E�^��=�}����)M�&�>��V����pc�}$����]�,k�O�f	��PHEz^��k�%|*����	ȗ>=:��4y��9m3$��+P�tH��0��F73ڕvB��r�nZ�Z�?A�R�۞��~-ׇ�����hQ���/D���F������c �4����A���a��*"m����,���r��3~K��t��IZ�.�^�5�d�r�y�U<�cx�-!�����³���/��ll���[�;ރ+�����/���h������/��+S��u��8���|��vNS�����e�K\	^��]Dq+�m�A-�3�1�8��H�hd�����'�cRIW��w��&�������Kb?�^M�5mO_�?Ś��'������I۪�������<��惋�J�
����^�J�q�[�Ŵr��B��[al�r��Wv���ۧ(sי)��?~��M�#�U��ik�*W��_^+U� b�F�#`�n�s,Oy�ӽ�����r�K�"ZAʼ��9(z��� �!}TQһ�K��n��E��e�@�y:W�������~��{v����n�����Xyϻ�3�� f�.�um'��ٿw�����7���Q���UZ��߰�������b���c�#qt�
�~�&�u�&�4b%���u}ǣ��:��s4���Q���ٮ� �1y�+�s���[�<��Y�Y)�Zc����*�᠙��� �:z��N�;��Ңc��ID��Ƿ��7Iy܎h�7�~�7GT�B�q��D����z|)��<_��O~{|٘�!e޽��KB��9�*�_�'���.�|�d�NԺe��0Ns51���S׹���ϫar��
�T��h
��h�l�i���y��4q�8w
^6��o+#����w����V}Z�	k���v���Z4m#���+=e�������̪#�#���/��|}ص�4�x<�G��
T$|f�s�z�2M	���t�����%�����Qҧ�A���MQmJ֣E~jаF,�;��nq?H��K�f��#k���.��E�G�p��ǿS̢�}��4�=�%��9�'�sEm7&�n�MP)���M�nF��p )/�(~h�k��*����FP�-h��B^D�!��ɧ�k���� e���l�A٩�7B���a�N��_�Ub�f��l� ��Oo�\��v>*��h��.��>?"�܄�b��y[�p�����Q|�(_��7����3�=�?�iy��zo`�i�Ik��:1��h���Db��G���8�_��nΐ%���q���������p����:� S����L�ó��$�?����hkϻ�x�󬭷KG /���U�M�L��q�8j��EHv������k%��X�>N��@[L�fRB�J�K"8��qM�*Mx�����mܫ1i�a#�i���[T҃��;z�o��j!)K���1��f��;���U��t�>	�Ed!�i�U�����VR���aV�$2�@8��+}#]u�-]n�����Y��!O�G�)o�����v���p���&o��[�a?ҭ�q�1����9���N�5ѵ��C��6�Y>`��~-�[Qn En�O�[&��I�!���*���&f��?k";��Os�Wr�x�/���DL��7uC�!�2�yLa���pNU���E0ϛ��T�޿�*��>��-x�`\�}������qN�x��	,��ߧ=	�L�E��u�p��-^t�Mw��f����ز�]���_G����"�E�C�Δ��7Oã��+�J��?�[�K�Y�4���xp��ٗ��[a���R#��xB�/R����I�/���L�Oa���&~ ��j Y��C_�HH��N����2b�$�oV �*3��s`�Ê�C�UW�7,�x�=��!���?���jzlx��L*ZK
�+��bv.GZ�-F��Qg�e	�oƧ+��+[b#�(�C}H���6K�)*'�gb4���CA��q�\%Pj��TE�ol�����D��(�����h������i��� �m����14QV��Ens�����à�v|ﮠ�����G1�����+�������}u5��K���ٛ��n�����&�ؓ�odu�&��2�H��%��� �!�p�.:kѰ�ܨY%�u{�3��̰e1Itl��3��k?��MTa0���. Z�n����U���p�T�=����W
Z>
�	�#�o����;-8��=��&D�(O����V�� ���ϡ��E�I$��1���CEIt�z� a�r���H�F��5br��.����Q?���
�Ec��:�<�"R�zC5Um�p�Cd-��o
��7;��k9~����6�����փ�]��r�C�`\ �'����`t%ߟXV�kUU'^-u�ΝOi�n��Yx����\DT
�dn�U�,�X��]s�FN��$��!`�;�q-➛s����_�w���mMF��տ~R�ߠ �ˊi,$��U�N����K��B�c>]  �V��E�E#�l����_��i�&�΅�8�!06��Qt������>����M��C9-�ZY2����6]��m �*������bh����,��>'�Oz���z�$�'�"��ʣͰ�:�T�r	%8�Z���ZS�W9t}��LU�k>[s��{���|Sl?7���6�xH���cS�/���6�!����<�@����©z4.�K�����"/M�.Eᵪ����L�f�V��1����$t���rr���s���1y��'�dG�Wܿ�3�ض��b�A�jn�Y
kZ�df��p�5�6���;�fɋ�>��u�x3!��d7���)uրן�kg*�����(贵�v_�p�`�s/mg�z/�WUG�[�h4�MPh�D܀�{P�7!_��O��^�?O�W'ְD�wa��u���rvy(���y���HpbV4����ן&?G߬�a�@�&e�`�W�IG�1�u)��1��,�S
�^��`+^��%i�St�<ɸ`Pe\��|Q��7p��d hj�wi?��i��@(���y�0����g�x�5�\��V12�_�Fl,svw���D�_	�s�T�"�����7%�T�VS��v�U1�e���ϝ�Z��5+�Q�01����Z�8�H��BV�I��^��M��?�K�;��Nψ� �y���6�F����p��ʜ��-�\�
R�_��b��aퟣE��d%����q0H,~�p��K,���h�ݠ�(��A�o:N\`�8��W�Z��~����՝}�yk���(a	���@�_�7�	��g;���L՜�5es����E�6?��$S��`TwIS����GW<ϗR}ő ��L&��Y�T��4���Px}�� ��,�t�����#�o!ms``����հ�Ͳ���p�u��w�2��E��I��JL�Y��g�k����K8&����H� � ok/��,X�d���M:�(|�b׏z-�WЉ�Z;��!��T��p�DqHh���Y~c��>�r�<y��r���=�}�b?�qd�YJ�n�i�x4����U�6+T�B����_�6���/����r�#�Ut#>mWOӹg7☨6�=���"���3 ĕ����s�c�}I�N�PǞ�}��Gz�� w��1�r���H+�<�,�����kP%T|��g� ��}���bfj�{�D�$}�>�7?��=V�b:�g[�h���Y*�)@�=�exr*�څx0N�7t�j:��VH�; �│���m[�_xx��sN3b�t���$�K�Y��D���p�E[�G;zJ��@��ӌ��mZF�-�/�g�X�M��Dԯ߶���z�7?;j���N��}��as��p�^>,a8�-MX�ڲQ�,��S�:�O.U�<��p���̔\!p�C���wZg����AQ�n���Ǣ��."@��o�]�t)*�p�]ғe�.-i��?%�m����5`�!��i�F2xv{��%	��M���Aū�����3q*��e�|cl1��\��]��I�x��y�w��K��H��9�m���1�r�B��:���p!b�}-�"~b3e�����C C_
�g��/�~�i���$B�1� �M<}IsP5 � cb��7V8���׸~��g?<��^A���V�/B*��V��}�q�MyIc0À�<UD56��/-ͻF�y<��n ��HI���֙��o��z4�ᵢ�y�����)��O�p��������ǜ�����9bb�7�2���׮��!��v��J���5`�$�m��L��H��������������,Hxri�u}f1��Y����0v��z������J��9����)�%t��;�J�=w�&*�G�&���9�e���I�"�)z���y�M6�I���)�+�RI��]|QF-�rjB锗W�n�TL5_1�����9mUf`P�;=��  �D��E!�w����v����W���Cf�e"�æRV> M
���8���7 �w!���O��gFw(ߠ����5f�je �O���^�u~:ףj}����ĤR�.���4�U�s8oa�̀�zѡZ(�4�i(�_*
ܳBaAl��3�3������wP&
YV	9������M�D$0w�A5N�r}�f������zj�08QWr/D�+y�/J�����>�(	=.��puMC�d��F�=�W��v�(
�������Ks�$jj�%����bt��х�/�.Xq"��AT m�,�T6'n<|n��m��$`�S���==�ᆮJؠ݄�3ѹ��ܫ P�ֳ��BSK������<��κ{.�o�����g��O�yb;!QWt/d*T~ܽ>�8{>c���WD��h
�����&������*�����'���?pd�$�:T�\�g�YD�Z;ՕO�ȹw�k>L��&�}A9��L�	 B>:CǱ��� �
��C\�v�n��t�v5�d��OKW_x�����A5������5���YR�e�ʘ�=Y��C�|��9�d���`���Nm��Z�ݎN�H�I���C���ߋ����A�F7\/E�yB�O��p�̽e�"�٭/6	�
1{��\-�1*�w�^�ۚ���k3��]�)|U���Kڐ�G���u^�2CQar�c��?:�����X�`�՗�
������8�x�]Jl���:˜3�ޯ��]��ٽ/.�/��EWD�>O�<@Ά41��5����ݹ�-+W������.��'��>&��}V�,y�'��bDO
\L�C�D���2N�CC�� �����C%���H�X��C��7/���ߌy�ZN�͈�c3�����[����d�h��Pt��jD���>&��ϢYY]^@�}��2��"�Ί��)���O7{n�d�K�����Ј�D�B�q{A7���'�� ����s�$T�;���PR[��ş/�y�Er0�x[(MY@�"�"`��YF%6�+3L(4:*����J������o�������n���?��כk-�u�_�G�@�:r��K��F��z#A
)?,�I���&��.�t̐&U?��%��3f���1fCI��^��|���C�e2o��t8��Q�s�~���d�"NrA�8�M��䷲�T��@�ϟ�١ �M�?�H} �z �g`��)���5�H��Q�o\�o4���B ��fr}���p�޹D���@�;�:Kb5�tُ/���ۯ!؀P����G������b��.)�K�u|k�U]A�+��iv�b��h0P�L�@�|�61�'���f���R�|\h���]�BޑI�0�EԷ4�'ߞ6=��zPti|��rkF�N�����W!x��00Z�KX�x�|��N �F�#7��Bt�ܔ�<�U���U�E�_/~��mvz�Uiw����µ��XnnD�+w��f��������]]��鱬����"��j�q"����Z�hd�5��\�#�#��ƿ�q�+*��D���.>�W7��Ð�,�k�JNdu�3�S�*=���U�i��ߠ�q����2e�K����^c��f��c[�I�w��ã��њ�j5+�p�@�c��'���ȱ�hӑ	W�X�\p
:4DQQ[��F�J�A(ʴ㡫`�`�;h�f�UZ�Cg6.m�m�ͧ3>�ٱL��l����/W�;Wapi"N	�l]p<e�!�堖bwa�ݓ9'AA$`i�ﺦ���o�v�L����Aet����|��+���Ԟ�4yyEӡ�l��6�Ax�OJ,&�6�z����	26�3G�Y���NRB~�iv�z��u��}+)n�CݓaDMu�Q�~%ᢣ��D��%}���ee���&V�}�?n� �*�/�N$�T���i+�\,�J�H�.2f�XO~�L�"	^�p�J���B�L�+�����w�O/����̎R]cF�N���}�2HT���8��x�g���:}�0���"�jͿ��˶���M���%�n{]�<$B��<�KK>�f)�Y�*��]Ӹ8��L�F��|,^�'��i0Y��a����ُ
z*i��-�a-���n���6�|���fa����C@f������Z�I�#���<����ebK�+�E��ؿ ��%�4e��[~����p)c��d>�s���l�mZ@ �)K�(:1 �%�%*���M0�4:����~�;b׍G�@��Q�us%��7�ಪ��y;?�8���>žk��>K4�~,��>���Y�ε��y ����"\�A�K�Y��r簾T"�D�d�+����?)
�T�����Y5�}��MY`^D&p�UW�_%�J8�ַ6��Xھ�#"� �:1�L>�#~QRs{�h��T�wXQֵ�@���ܰ��E�<�������r��Xdۦ�/��Q�o+3푆j��7�U�ZcΕ1y�@��i5��B���h�̂c�Qr������ձHE�X?�=S��F���;n�N�@2��Y ����o�\���8�qTzeׂ���uu?e�O�F;��Pz\-l�JQ��7� �O&1n��I���/~�z�bu��玛^�	B�W�(Hрa7&Z������k��?�c����؜x��C=c����|�	�l���ˬ�kCE��3�`ڼ,��/�}��iU��p�.���-�����z
���n�^������n�.��n�����.��CBi��w�����}����9s���;s߲y��X>��ȿط��ю���s�e����\�,T��P(e�T�ރ�Ŧ6��#���1H������Ħ���e���u����	�S��Qj��*�	�7��m�Ɠ�H�ե��^u\\IBhh�$(-�Aȵ�f�Q0$0Lu�J[Gb���e�(���Y�OX(wMy���C�FQ���<\j�ޫ�
������#��g9uM�2P\�7�$���l���&8��a%Ұ9G\i!���1��4=8<M��D�sG�R.$8�t�i��?O		���{�)5�A��!i!�+|cw
W(+:d~h���'̵���X����8)�]�H,��f9C�%�c�z���CF��"V���ĊەC~�E"�Q���j�Mi�B
����ZS1j
vn����&��YHL��y�H�R�#�5�������a��8�߉���l�~�+�YT�w�?�`��;�-�[ڨ�=��[H����M��	e<p�J���I\�V�T�IN��+�G�NPʏ3�_�6��ް��&�C��4����l�;�)$�@\=z�,x70�{�d�|��즨�<lyg�D�ж�����gBi%����&4t/��-�NH��i�~?���y����.�b&��Y]T W5���B{�zGL	���`T���{����F�Wخ�9{��Ӻ���t���|���{v�e��$M�4 }d$J3v#Bxn�C�i �pG�����p)���{��3a�_���.�|]T��5
*�I�{���@��!fo��p���>���l�C�_�Ptq�P�D�Y�`�a�Du��s�����8T� ��:�	h�����\> ��/P��l�xh��s�W.L��ў�j���ޕ_m��6���+Wb=�ڰ�l_,*u3��W��C��Ζ�q�:�M��W�c��\�>�	��q��H+N��7C&
�NR�Y�������()������
ҍ�� � X)����&#^����Azr_2��_M��!_�a>ሃ��k>������Q�Im	�imD�v.��:H/�Ɠ~�m�7�Ó�$�%��Y�o���(l����p�Ψ�1m1�����n�oG��$$�aK����&�ew�o3x���ʊ��FGX�:��2�(l�j���p�1C���4�&�P+�eZ6:{�vpw8�pD�
#���P�SQJx�����G���q���͓^�3��Eo,���s�Ϩ� K�&9J�04���yJ�h-�v@���P�����TCoͨr8��%�T��c�_W�Uz`���o����O6HW�+��Н/}!��7��5h���{ 7�'E?�v�F/���K���A�ra���(a�$fx`�ġӨ�C����Of~�䄧�DG�
�R��?i����p-u���G�C�"��/6�u�X�A��\�	����  ^����-��	T�v��
_p4�<yk3a�7ü2͜��:��섕�Ge�"�l���8"w2N��|�yb��e������g���2~�6αv?k1�~<�������ƀw#6�[�E� ��F��F �Eڂ=B�@���_p��\��^�ƫ�zDǺ!�fK"�\�^��/7e�vA��WzD�,:\�����C_#jk��F#	T�QX����汃H�̉�i��2�-��n�����%��<�����O�9+a�w'�߿G�Fي�%MH�_�:��*��UT�ڄn���Ʀ�e�x�LD0�?�E�����&��5����#zf1bqf�ۥC3�-v$/۷�ùW�~wbz�^��Y�~���|#���FX����oɺ��PYH��O��6��|���6�	�DnVW��!>"^��m�9/Xg��τ&d��*��FKD��G�Y�g��#E"� ����� �#Vٓ �=�{�h �����B~��GL�1�
����*& {��@ 4��B�����:%1�`���x!�	��k�~��:���,� �M��(B�������q
0�����c���]��L�ڈ�L3! � �7��׌��ЁvY��x���7G�$��dX�@����Ƙ���]	���2�C1�\ ى��i`僀|	��(`���`,����� ��kC`?���<��_�=��8 >��?rQ �HC�9�L�_3�L4���杋�� ���@�=���SDv1v2���Ձ��F��y���|��}�O���c�ՁG�z����{>LsMD8<D7�L7(ژ�<p%�,7���p�D����fi�@֩�7��\rB�;8�J���R��U6ǇX�6M��T��&����da\�PO�#A|A�A�m�Z};�$��	���Y�;�}J�O&gI�r%���yB$۷."�X�(�c]0�(v�"�3be�1��u\����P��T��$�Y����xu���(�ڍ,sM���X�b*>O�qGv 8x[PR]��f\�`)Pg��6���el�a�򠗭��Z�(*����g{*v�ct���$y�"Ui1j����H�"���zH�'���td��oHL�#䃴9��^&@9��~쿏�NC��RG=��Y8����$�@@��m�T���%0� ���$G�^0w+aC�#$������ט`�g$�L���Ag�t۱��06��^�����֩\�0�G���R��)ZfΘC�<(��}Z20���8��i	�9�ؖY �m�����7�~Z��x��ե
s42w��B&	��J�Y8�ޙ��:��F/nǬ�2~��ᩰ5�d50�Ӥ�2���S��W�d�zش_ْW�@�����9��Yz���G�T�ғuhm�a��+�6���wB��9����20
�A�� M]����Fa�X
@�~0I�{<�۴���)��|��-X��n,���߯�0	T�4i:���)Af�{��#�LZW���;�����z�;�K�Z��y�p��R��A�1O��GK���ɹ[ۨ��%eZX.�n%+D
O<�\��F ���?�'AKIɏ]Ϟ�w	�ƢN<Uj$�����F�C���������U2e�T"���5��+Čp��y@�k\<l!�mt����_[Y�c�Ld���B��RvN����Ǒ��m{��lbIJ��&�8�\j�2���	�|��R^0��B�'�JBNG���(�.���ç_��L <� ��b�R!qh_��yD��4)!�s�(����W�G������eպ��/<\
����,.$��W���
��ݍ�rI�u���c�Tn���4�����*7�]"�W�%ͳz�������gZE��� �P�&->B%��Q����Į����9�x��=�r�:��7��M��w*	�ˑ�g5R�uEy��tk��)���%�ؾ�˘�yғX�\+��Y��? ���N0
�)f~QH���.�	bs�_��Z��2�5ս7���V��výNr�Z��h}@S���ߋNe�q�6X?NmT����m��m����ѹ��_#�v�$�U� ��~��j_��H�\0��@��"<li��ț�l�n���AZ�QRJJy$�9F��Ht,�����H���o5��kfb���2W�'x��;�1=?�0�KN��+�����c��;sXWQ	G�"��4c�����
A�,۲خ߳W�9�Uq�W;s*�XA�,v�_M��i�2�_�/�[7��v�HKKW�yy�|Kx�+Ǿdm>�k�_��z�1�D�*Ll5�>C�Q=�"�D�emP.�X��]����qǥN�<��ieE��J^ş����vn��iU��}�g|�'�ڴ��	��\��KP= ���~�Hy���1om=��$V�㝟x�t��^b�a��&(Q;3�5X��6�d_���ǣ��S������a����@��գ�n���ބ�adm�#�|��PmP�n�f��T����TXu�y�u�U����_�&ݾ~r��\Y[/�~����Uj��ū<X&|k@6���3 v�ga�[O�xz���F��3����?�2���/��u�O%W�?������0ޫ�*A�u0>�H�1ޛ�%���OnS�qMfHH�(�$�k��w2��+��7��CDȤW'5�\���ޛ����ʩUg�įo`a�F1{�r���R�
���!O2���]�v�� ;�h���꣞��ХAX����5C��q�l(��8���j��6%@� �E�US5��M�R���	�]�]0���G9q�����)�=��G��C'��N��"�[�I�A?O%֭���2Н�����糍�_YPy����v|~7�Bf����,֯_�q�|��>�Lxh��l��Pm�,��Hx'}��W\|��r�=u������:*��<5}��Z=�;O���/�:��KU��g[���7\k$�o3e��X�_�(�\MS4�q����usg��M�nGG���%x7-_�]�O�U�Zĉ���v�X�Y4��-����@�Iŧ���w��o�Ec~�'�6V�E�wE+t[�P�##qJhj��^Sm��>�i�_�e���U���J�v���F;��%�����M겧�|���3��Mh��r65���v�g��4�4���vn��kIs���'噿�t�1�=�����2�xj�ٶѲ�M}@�L�+��	6�5�-c�f.m��f{��}F���'�򢜹r����z�F�~[��������g,U6'��S�H��l��Vos����%G$�6eH|�{{ζ(9qT�H�R]�i��b��YAަ����lXϤ�2I�NѶ���QӷQ�*:���n������0F2?��>�>�!��ԿY�Q����j��3I����֑����	_��댏���5�Ŧ�ٰ��f�@��j3�|͕���rX�0�3��������Z��*o�J��i������Pi��C9j�(8z��hT4-�J'%��O�,l�;��]�`�f�()�;�f��l]��������@j5�U8�w֢���}ޡ�<~H�	�T8]]�4|�1x[�ت�fp��
����m%(͌�R�vxr����_P�!+M�5k1��s���Ό�4���EcK�Ϙ����ٸ��R��>�m���6:б$�Z�� �Rz��7�v͍��8��p�]f�}wδ,F��@��T(^}�;�/q�j�O䝮�+���`�&��D�0*m՝�E�+4f=zH�\�,1e΢qG���st~^	C1�;�q���'������e#[��ơ�w�J֩�����m�p�Y�~Z�¢��O�5*�Ҷi���b�39n��\��]2!�I"��g��q�����?Ȉ Y���&�/q[1���ϣfM7��>=%�w����]����x�5d�`�3�AtC���﫷kMM�hGɑ,z�2W�辣>��!�^��*�[���&
A2�z}[HM�]�I��������h��ao��|��՛��aC�F8�����dɈ�
u=ej]&!/��I�~j~ɬ�m,�f�B�̇�8ң��Y�6<��7/�ۭZ��v`Nc�����yQ��Q`@�ڵ~G
���e,a����O���2����D�*��4���,Xw�z#_�s���ڝ��v��;=�ӶF6��-��ua+C_�� j�'6[�z���S����~�M�'���cg�Cxwoh��P���x�&S��U�\��7��Ļ�����6{��q,%�Z)���j�C1�y��&��T��&	�M��F^�r;m%��jg�O�@��D�8^7]�~�¯�������_}f]�����)XF�p�U-V+.�d�U���6�{L�WC����8��N���w;t�v�m>��s��WV�|�>�y�m�N��Hr�1��߫9`�S���U�d#��C6d25�a���`禡Jq�[��T�f�;��]WǨi���+�a��ɡ�'YY8)c����r�R�ۉyh����=���_o3bͻ�KI�#��ݿ�g����?�Y��t.n����N���0n��[\G����UC�ۄ� ���z�".&,N�"�2&%K�ޖ���G��p\O�g��흴׾�E�@�<R�վ���Iemd[�������mY1,y&<Q�{%l|�t��V����G��F����5�l7����H�7�J�GsӶC���lDkd�q��y_@���T���?b������g1D�~��6Xq�vV5�aI΃���c�������C�d��n�n➦��n�Wn�K��;���^���ܤ�9�㜏}qK.��y������x��b��j
���J�Y	����[�ͭ�2�>�BR�)��Kҋv���B$����I�k��� %����?�qЕ���^'YӘӾ�@e�KN?�#]���ڨ��R��'����ϵL��f���J�7����ܙ�Ÿ� wL�P�7� �{��C$
yLGP��1 }��

ڈF� �/
5�Y����R�j��
���EI��;��x�'̵�xO�W_5��@�K��ymn������z&ju���-�/�Y�<|TK�3.7J���Ê�Y�$���UJ������]���ى�Q�I�+�1��o�I�p�rz�Dj�n߁�����RPk��ت'x�+�\���fo�gG������[vxʴ�O�Jc��!΃��Eu����K�ndUrR�
��Y����C�h�#����樓c��ܻ�@R��%pzn/Fܶ����=�=7��� ���!�����dU��s#�=�aA�~�הå���
��_�9'�TM��vfڲH�#���\ҶŲ��gB ������
�XP�[I>����]�E~�v����;�315)�YY�R�C���x��?���a�Μ�Z����go`��TЦ"E;c}k����p��A��5�1�Q!�Di�B�u�op�8}��=^����uO*�����{.���8��$+��{?[�]��s톇o%L�ޔW��P��"a�����)-�B���]l��V|Lq�{⟤�g��V~+>=���o6:4��t
��T(������[��R{R�8��ɻ�5OZ�8f�r��7��d�W��xb�H,4���84]��ܷ�䐃!�=;�����	^o�FL�#�5xE��x!����m������]�����IGo���s���%���n�*z�F������qo��NDG� 1BG<z�skA)N���i/%�oy����:ُf�Q�׿���2Jw��m[���J>��uD9l�F��X�ٸD���I�)j�D����C��#!�_������zؖ��HB�*Z>{��9È=��A��8/j�jc�؝���H����c��,��P���A��g��j�v��
)�l,�����+&(h~��~w�����:X\�J|�$���N�l���d*�����9iV�$q�i�⓪9)�&ڵ��9�	�ߖ+�,�4�J�4,�^��u��sf~!��o{54�ƣ�dMv>�R�$�����a�@~3�A#g�Ol-�l�~�R�Xe�3I�x���s����@�M�\8�(�:���&hH������X��<��PR*`���ӧ({ *|;S�H�H#�X�7�	_ ���mS)�-�m��āg���b�"k���g��3㧣S0�m��j8���F��~Z�h�Ż���fC��3�ë�E�$���������fo.+�'s#�ȉΥ�Ѳ#�%n9���X����2#�S�O����s=�|�j���7q&$�F��6�����w�8(�;�e���e�Z���@�r)�oo�Mrko7�g�Na����_��!�G~7��{��F(�\��or�|��z�p�Ug�T��Pdq�ט˲��e�����u~��Q��ޫ{w�G|��@w�
8L��x�����B���Ƿ�͹Zt��mu�+�_6����eĄT�4��Y(�YNpHX0�\��d��N��\��"��qk�b�n������ڈ�x����/Ls�z4"x��_�Y��D�n����aj��.����Gb��(����L�["�v��c���G��K6��!H�*FIs�������������W��Dl��1 DT�����L��z�T��=_K<,Fg�e ��
�d�td3���y���W&��|��0����o���9�YǙ�fC�ȇ��-�Û"P��NG+�O�\�u�O-@*�r�v�"�⃃;de>r�k��q�i1��jI[W���(b��xE�Zf��l�g�??;zFR��'n��pt�y�z�O��=k�AGl�U)���]'X���8Q_0}g��%����n?��:c��$Fw{X���{��یVDn���)fw�>�]��;��3��Z؝W�.��I�OɋB��M	�u��:ݖ����:.��!�MBP�]P;DI��y�ʫA؛�!I�G(*��4�ȷ�2nn6�P��P����堁Gp"&f�E� �������oE��g��9U����0�����������%� �i�ȕ� dR�p0<U�/Oi���P41�����5�7[���SL©7k؀ur��Vq��h�����e���,'C$�
�qC�?>m�T�)�`
��P���fٽMsa�Y��Fq/p��Q�չ�\P�I7�@�!�#�,�Z������|�BZ�r�M}�FΞ��{Td'��!�ԙҝk!�j3��>8Q�	Bw�nq����#��v��yjpؑq �h$]/ �L	�RЛ�M���]a�c�766��-Q��#$�]Ӳ�כ���:��O�D�*=���(lU-Z��f��P�:#����6���
����w�Y�W�f������Ê��8 ��5�ݜ[���~y�&q��  ��m�P��q�R~&��/�p ��/Z�����]�4�Q�TD. ?��~jU_ۚe�gi��ݮ�Z$j�hh`~��rkG�4d�	�)n
���-��모 �w�t�r&�gqo��<�p0d��q�S��i!��g@��	/~ՓRٺ�����f���fz��$л�m�
���|�9Aշ���OO�7�O;/&�NO'��[�c��j�����ȧJ͆�Y݌iU���:WR%^����`t?����vW���@�9{׀ϥ7����~�r؛w9L$h�C���.G�Զ��翃8�t��WT��;���ά昖�Q�a�4Й?K��lji���&�vS8`��$]�^�������/�k��}Mޯ�+�}}x`6�y��]��śY�L���
y�b�4H"=wL#yq��-�����zI�����w��)j(`^%^YM�;��k?H�#`�h^ȴ��z�Q�mL6�!�ޮ�x�6���~5���n�o�>���d-WQ��@?��[��2ş�o.��c�vB�J�k���Q����g�����3Y ��&��!���+�¦⽑1!C�2�؈ٿH!�ԄQ�Q�)���&t$�q;\�Hrl�B��\��J}X�B%2�>�H.^�������M�ڃ��Pb�2��V�ـ��fYԆ�u�]�냮C"B���N�8Q�!iTu)
r�1�Ȃ���%���`�"��V��}YP�H.�ʗ��7R?�=Φ�����^~)@���)�i��	H��moy�;aW�Ν�l@�t��`H�����5�����"2$�']JE�!�c]�.���zs,ܷ-��(X�nr��+ Y��A�M MQ0�6xYM���r�5���7�3�Pfn�=��T��y1��.�7��d�:@�{h|������8O���g#ٟ]�╡&;�x�v�-���[��)��B��gRj_ޜ�i�^!/-`	���h�вe�j��J&A���3XE��%Ƈal@��H8�6��t�YJ����Y��b�f(���,{�ό�t�)���x���:�����y-�%cz��n/2J
��2���l���4�g���$�,���a�J�G���Mޔui\f�����������?�a�����97&gi:Z=՜#��
_��]�;m��ځ�[����_�V�$.k� r?����srw8���ڲb^㊚tɋ�� ��qj�^l�yڒ���>��P:J���Yo�l�?��}1^�f�s�����;��w�� �W��*��W����ï`���m�C�����j�-_�?԰a9��@������N��i#ˁӄ�.��l[�g�^��:�n/���$έ�(hJ6n��؈��v�5a}��&"�g��9Q������)N��y#��:�y���Ȫ�����z��{����fUT���l�����:���獉x�{L�ʴ�d̔��On�c���Z7���s��N��r�	��Yǆ7�pȟP�o��-S�Y��>
���Y����& w�5�Z�~qI6|�6ے��ъR'f�1�ϊB�~R}�v!3�����N�?_o|xIm
p�0!��$���	�g�\0@S(L���1	�s�{�`B��-��^�s5��GK��f�Am���+>�?{\�d:����ل}�78�E�X<B�H�U����0yE@JJZ�٬�#�̌�M���(����P������yO��y��oK�l��2�˦5�"��b�L� ���ojh�uk߭fu�Ƣ�4������J�U�k�珙�Z��M�\Q�z-6D���za�:��W�>���N�8�_a�[�����uhE�d����m �q6-��P����'�F>1m/���?���;�b�i�fy�ۀ������^�(f�� ��{��n2������0%ox]�̙�]�ޏg��`�yv�O��~�̟k��@�|�z�.9����2���U�w버�vۚF����q������+j7+Q�-`=<�:q����7�SXpd>>�H>n�Ds�
��*�}inv=�GVB~x�I�K5L��,(e�%Ԓ`X7W�*�x���ԗ�`G^���u�J�Ro�Y�H*�.�")��k�۽Wm��Z���/�vI���-o��4���ޛ��_W2Rn�E��� ��sv�����/^E-��rȅ\��4V�s���u$�q���>~���8z�[hr2V�E�]�U��N�l��癭$��c-v�R�/���Uhl��y)bxnW�n��e.���`��L@���{'���+�T��zye���:�LT�J\��]^6�&D5��
q��?*�w�R4�WmY�o��oߟ���A� �n����M^�-���7nhw!u��
�4��7"���V{x�u�����#B����1c��G�e���+�\���!�8�.�˨�����d��֦,�j��j��>d|��1�$�T������b6����k�(u0,(�/	�MB��N����T3���h�u�CB�g�˞9�B�'K��l9N�$�M����b������Z�ga���*��b�HH��4��@gͧ�ݏ��n^Ϋ$�%~��U�Ȁ�����X�4�i6?B(��Zu�8��Rw��'#��߆�L��Y�i�閍;QR�6s|�)́9$� ��B��q<_��#��|a\�#����Q	\$N��=j^����H��z�Mrˀ�y�Z�V�C��QeU�2�Sz���#"���s��i�2;�e�w��e�^��">�8h�62�̅�%X�?޼�V��Q�=]i��]o�=�S�gI�/c�oX�q"Ǻ�mr.�/�rq���>�s�ػ[9�_���)[m�rg^bURiE�Km)r�S�Jn�9f:*!2HÆyf�N�S8�X;��j�)]e�S��Hz���g�[^t�#X�tq�9�Y�q�p�s�����U��y��J2�n`j����c5e"�"�n`����>�R�����\��tg-&QՋ�6��V|����������t�b4Z�f���$�����"<8���8E�$���0�l�mڧ�#|b�*>qV/�����f����J�u���.�����D�<�7$�D��<��t6�+���T�9�8�6�'�������"�f�ń|ؿ�,ȷz'�Ũ��3#�����k"��b�%���xN����n��-�lL��&�[fg)Q��K�4tBc�ִ���{B,��5O���͟��X�6��U�-�����<������ރ,m��I4(�GX����󡤊d�-t�8&
W�o�M�y΂B_Ү��.dYZSd���d�׵����rF(3o7�����WS��x���O/˚X��ұ3�����TA��B�u�?��>�]��(0$�y:l>�	*(���v�a�t$�v}B� ��x�!�v�΀��Nm�w�7�={�}���v�n�m�	�#r#�y��`P���}&���Ԭ/����u!,HRlX?�y�h|��\�h�1�w�֍!EAN"uv���]��C�y��$r�~0z:G���<nD���|n$�CՋ�&�r�Nԝ���8��yP4��<A�❎_W苾��7��Ⱦ�����?c���gz|j���ɲ����!D�d-���.�hF��x7�󡯹GJ84uF�ɥM)Lbj�-!�B�ǈ��8V�ܿ��%3���=6�O��x3�⵿D��ў/�1�Agd�EDm�8�f�/�޾����OE5��o�}�adv�ԗ�斾��'�D�v�VɴH�"��"-��s�kܘ~x����X�#�"}d.Y�;Dx󼤕m�-�_�n�GK��x��������߶��&H�{{�4�k�j4�pr�Է�-A��>����{������oÜ���x�G��2c1����p��4�]Ь����`��]T���z��~�fQg�(e�x6�M��I�=hgH(�]�'�?f���=.�[�H�g��/�h�)�,�|1I�6�d	L��!�zt�������@��Mh��ʟc��ҵ�m[�s�SH����|��f� q�d�pU�~�w�r����w3�e��YI��R�r�=ٱDH���kC��Fl��y�w���3]���B`M�����h���#�E��H������n8��`퐲
�K�n�EU��5ii\0�$��%�Md��Ekl���!<�E��1��[޻�iB�)�e�t�}�������{S�@��0��0�d�yQj�S���䟃01��m�K��U)\sB��ŦMxBG0�1
H���&J	>�q�f[P�f1���@1QrX��2����գ��Q��O�D���s\���L!j5'�Y�D`����g� �0�8l;��
"��96�)�A�x2d:)Da��R�,c�{Q���JJJ�@�',E�$��̚$P�c��t�^��T�2�%%���c �B�sCxE7�?1������YD#PL���|���>���͠% ��'�GH!z$A��_�L \F��@q	�Å��B��,���i$�OC�� ��A l��DY��� ��1dL=v�)UȘ�a�7�Gm�cF�멂B�2&��y���<d��;��� hMA�cԐ��@O~@$���(�_ � # �2?��	� \ ��Lq�z�\l���	��-�ƀ���`˷@hH���ɮ�TK A����_�V����d���qBHH�����^�
Ї�	�U�7��� �4B�O|e���} nVA�G]".7B�&� n8E�`��-NY��9�"ȍR�jV�Y�X04�/
w�B0��C���� W��}k}���G.LKu������J��ݚJZ����\�Aue�\D;j���ҍ�n,}�He��
�su]P�����R�֒�y�z����K4D; f�hp2f�U���n�J(��t���!�ȡ�ЬGXE���a<��|>kŏW���%�Wt 8Z�� =J"�%�ݖe
�֢ʐ������@�]��z�p�}�9W�<�II{���eL�:p�)�Yc�z�)o8�PL+顇���>�ô���j���������3<�0�1X�#=��q� <���ML+�����a����ĢD�oH��F���u=���@�A���ւ�B%����p��С�N_��Q��ç~���MAe)z\H�T�Ѫ�|W��LA�2h�ܲAl0���;1�nO��%������z�0����RZ���C�d�Jf�O�[5�����.y� 0�̓������. u�OH���ej����#��J�<w��&%>X"њ�{��f�.�%A��H�׃5&$�2M�K���	M�
�#��Ats�Ε������=Е:�+�E�"D@�����YDm�����u�"}�~nyv�VZ1� �$�VLF&�2�R�6</�Ĺ��?�CaN'��}G�̈́����CH+�m�+�X�9����`��\I-���n�C?���B��p��s��Fɰ��'��������ԗ{��=��j�Ik��%3J�mw�]I�bO6���C�V��&B�� Z0��6{���|c$�4%l���=#�2	�9�F@]#,KQ4a��A�[�����x�;��Sk���䖂�Z�T5�u����[)"��2v��wA����[����?P`3J(㨈H%99Bz_��\����b�,�v"L?��D(L]$T��^H��0�a(�55�0����J�JN�8Jəz�!���Mͺ�Q�!۫u�4?�k�� F�%,���,	���/8})N�o2Wc�eպ��̷o�۪)�NK�wte������d����3��R@�i�:ޝ���z�TdrX��Z(�Bd��g��	���P޸=�:`�Y_0�!BOa��X��Hsr�z�)�u
,��(0/-)�v�z|�v��]d1�ߥg�i������ć�דɝ�
tb뜾�%�v���<����zT���PW}	�3�,�{hx/�=��$D�׼�<�z$"�Ӫ��.��`.����2�&���K���C���Nw�2�m�J+_n�%
dͽ��J�φ�)y1g�������:�m"�b'�L�pU҄���@���7��w8�� �0`P��(�����m,����>sl��;�ii�Hʭk�FKNr80ڜ3`�;{�E��s���i9��~^آ�GC9p�?�r7���#�
���I��K�i~[��4,�����0��`9}`���c���eE?�a9O#W�Y� =�f��с�-U������M��@��z�G������8���.F�?$ӿs�C�/��ԉ�6�j@�V[;�����	�A/(�O)/�B޻��+0'��u%8lG�`70vk}G
͂gi�%=��B^q<Yn�����'\Ee���םߴ�:�ۜ ������.C�^ڣ��k�tf�B���<s�n�W������ܻ[��n�͏c(�\푩{��]��zm�ٷ�6W��w{�y:���УPJJ. �����RV�g���У����̛�O�]CԳ"�vO��?���`�� �3=%I����@ޭ�D�uE&�����o\?W��=�ʳ���My�z��3����4K���g_ֿ=t��i��7��j��
v���������w��0����F�Ni9V�N�ibF7	��h�=[��~��M��z�tzZwv�����Q���dK�z(�l"`<p3�+�y2��_Z�����e�&j� �"�t�9W�\c�c���"��-�Xi�F��Vp_ֳ�\��rdL�r����;.��7�0S'�DO��E.
���EW���zsa\�����OnE��J�*#
�*8���B���DU�Ye�[Rum�FS�v;�Ы��
s۽�|�^��/�YIH+1]���5���Un'�+_/��U�	������|�K��rr��Vh1��VQ�f�D�Ƶo�6�x[︓�x��#"��5o����ѓ4��I�(�	lc�|&�����x���m�׹���c���S��8ΟK���{C�^iԹ��\a�����WN`��<|���&}��ix��(_}��*%}w�\ܳ��'X�J�h��R^�:�k�뼞�E����wk�ظU���x7��sy#�	]4.�V��t�G&�?0���㥿�7�;�8��R}<�(�&��;BMh(��A�K\Ҍ�x��B�:�5����d3Ld��U����w	^��H���>^v�v'i�}q"�sSl���Q�����t戻`��
+�����㺂��j��Dna�ͪ��D$Y�l�E�o(\&���a�\�?CJ���	+*��頱7�"~<|��:���o�'x�ƭ��ة���>?P�i�V��9��uP��ww5l ���6��"��1�r���Ź�����3�R��V��u}
��<&²(\@K�_L�>��2�I\wҶj�Ĺ�J
��#탡gSBjF�ƒ��
k���#���7�x�����FOQ���g
�?���:ck4��������Fz��o)�1;-;���*�[��?5 ���Mit\d���Ģ⇗�д��_<��+Q�ZQ64��Mւ��e�R��W�*���?^�^��DP�E",�̭.��u;���R�U��
?F�AVn4u?f�����^������>�P�_F���/��q�d�m�4�,��h��{qy�˾y�h�IP�?m~J|"y;p��$�R���F2�h���%��ػ�}����-EG� �E?��l�	���M�C��΄,yL��4�g���}��5�8�?C��.��p��٫4�mQW��,��
=	�һ6�e��H���x,g�:���.fs��@J�(���8\ǷĆT`h��n����t�w��f]��6��@�������$��,����}I,����j���66�P���k]{i�y�oI\��*&��Hd�O�Q�:&�D������7���YC(R���
Fwy���1=v4V�|˪����������i֋�Cpw'wנ	��N� ��[p]48�eC�8���w�9��StwuM�SO�T�HHĊ�IdE@H�Y,��[\�� ��o1�x�U�AxÜ$��i�݂V�%��SC�	"`t��e���9�D�x����!��F�d�������8smK�XWE����5Ua��i��Q��K�4���x��qS�Y�q󩡀�XP��Z�V>`]@}��Dx��D��v� ��l4P(po�o� �x�6ɁE�����{y�<jZ����mxR�-n����������*�rg��(��V�y^(<q���J��h��u[�,��V��ŗ_(=�hv�d���r����7�%0rW\�~��72jʱX�f� ����].*�m�2Э߉���s����:�����3��<W�#dsDX��⌬(Y}�[�6,xb�NM�%�̻첎���jyJ�]�2�iw��|l�hx�\�s�ò��b��45��9�*�p7ћ�yR��U衭��C��<&5_��)�	��x���rb���{s^�u��Y�ga�F�u[*Cr!�r��� h'tK��R*H��go�t��V�E�z�ѓF��=�7�w�R���o�UٌzL^�?��K��(n���;:�\i�4"t-�4x5֑_|��MX<�׿`Մ�}�G{"�r˶��������z��2q�^���?��f���|��G���Sr�s��&_����d�Z��2�_��]� &��w*Z�r%[s���a��(}�Z��gVF˦I��ܲ:���#�Z'>����dv�w�)��]��	�)tb�<+Րe�=�vվI���妎b���H�<v�7����/�z<:Q�?�q��M:]����u���ʴ�T��΅MR �<2v�/�J�@8��]D:�Q��%2gh�:}�,�i��9���o�/!�dwYV���^q�
�Ԋ-�m�&dl��r����뉤�*�U��6�b�M��]�y�1=�$�b����t�w��I��c�ȤR�C_�`_�ٖ�O�=yqa?޵��)�q��9����6X�|,ϸ�'0X2ϴ��H��2{�V���(��3$��s�*��/�q��#U?��@�ɋՃs�'C��/}�6���{��F�G�ۏ�\���i֡�Xb��{H����|���k%}�֝,7��`��-dI�-z'�8�:am���zE�Ǥ1�hڹ4'\7���+U^}�j�r��@*$����n$P�N�-�!p�ϩ®��l����r�Ѡ��r���@?�C�x�C{��v��K"��^G��N�WN݀�������51H�K��K�����e\i�NǺC o;�/�d�u����%/������(�r;��`���//���c�A1J��/n��P#."��h��~�H��"N4\veÆZl̘���!�� m�4,��K�j�G�iR!����۫=�'u�`'��&kt])mM�Fz��9��'W:�OB5?�����ƿ���ǘ��3.����������n*q|ij�fp�w#��*NC$�v��g�>�i�����_��<xT�t ��<K%�6��&�ƥ>FW�9 ѢЋ"�f�|Vwx�ơa�h��j����l`����[u5�<�R{3�-+������!�����)J/}���02.� �4���m��h��ލ���J�|Q�aw3�u�K���ɠ��\��կ� ّxPIG�PF�U�jd�,��rļ|��C?��í�צ�i��H����+p�џ̂�����#+T�
��N�z_���U/���#,��dQ��@��Kd��Ih��8�	��
��#w���2���H���x􍖟u�9BPCC4u����ۡ���B����1����n�{�Ȋ} �J ��L��eE�'RȖh"�/˙@owp�=��[��c]V����휾�V�R*���~��Y��S�]v��k;���e��*z��h�̞7�!&���X�Y^�	u��KP_�Y��0P�7@z��$�oC8���ғz&7RW=� �F|ƾ@�\>zq7q�J�b�dtՌ��](K�m/�����G!Z��U|�.�>��(}��~����
�)wp3H�2l��F����x>T�����5�<DJliYm�So�̭H�" ۦ:�j��t$�a���$V�Q'������|8���5���$����g����m���W3�XBlы;���O�庋�(C��H ���"�;�8������{ON�Y{��v�{�ͨ�
��P9)a �B"aO;%6ؾF�I���ʷ,�.s[��ǚBb2Q_�J �����[&���-�?=JP�/Z����o4��~_�(/����;b�L�U����I�ʝ"R�{"��d� �'ר��� �V���[e*W|P�eQ�ѩDve ��>=�!���m1��bd%R���a�����(�_ZI���?qб1E�d�.���Q��Z캨o�`NQ�NX���)A�l�w"H�Z���b��A�[��k���n�Z-��|4��
���,h��h3���&�j��|�������o��@Y�RqH�2葺�����}��`�c��-տ�Ge�n:�H����e��"�V�%J:J��B�=��i6�*"�7B�ą������6bg�6D��.��*rn��!��Х;bI!Գ�����B�X��jK3ʊ@���O,�)��/}(�7

��,�6�Za��Ҷ��7�E٭����k��Gm@\tZT�_���%F���┯��^%w�'��B���2�g�!�3���[Y5���a(1`��Ƕ��~`�uG�@���Q7!Ͻ���g"+z������F����I�?����T�P^B�G�A�W�����9����~��DcΩqB�O��z�w&:ss�d� ®z�t��3����Rm�ҽ��w�����nr��hy�"2B��Ӷ���ِtRR�mv�+�tY'�_=7L;�	vh��N��!��+�:X��'A���;���..�W(�j�5�Z1c��t��v�%�p�Ә�M��#��\@�|���/rW'��f�F,�[{�Ȳ�~���r����6Q�x윗�(�KPV�;TbJ�<$��jW�]X ֈ7�X��������,�R?N%C����E�`R
�܌���ju��	� �i�;Mo
V[�j�C��DS�@�+D �9�꿛�eN��n���q��_sI1�4+8����\��t
�x~��hyd���3�L�wE�l� S�1#q��"��������P�bd=���Q��;N1(�-�2_����b:
47��v[�;\��b�^��&�*;6]��{k^z�qл���]������{P��ǥ4)J�w܇�TS8&�ʴ����e*_O����4�N���΀%+�7z�)J��Y�ĨP �Q�X�����Y�7�c�\5d/�&9z_��b���	�of��p�O���O�9)�Id���1����(��{�ח#E��Of)F_.?���t�҅�c�"�t��{B�H�q�[�4+"#E��;���h�l-Ռ뚮��o�sM%ay�Q	�O_�~�oƄZ�
]!����!��[��z�*o�m�z����0��hL��V���_�yU9 D���ߧ�_�Ї׍���ޜL��Gα�[�>�˲o��HyC}�k}5��zuB!����rQ_�AR�wOY�26}�;�B�c)��������K,��0�3�̇���>�=��h��t�s�A����,	�u�<e"�l8��*����rP@�ظL*�y�X�,P}��mCF��^R�Y���x�j]��x>ˇ��wn%��l�ޛ�bq�4�[�����Z����~~*ri����{�7|�!�~�)�m~(���6��]�eHS�S� 4�-6�����V�E����.����5�+r��R~���1�9��lF�(Q�1��?��J� �IF�tJ�O�Jz�oO�ǡ�c7���r��P��B*��60�v��86��*`�J(�����T��y�S��@��y�m%As�i#��>��\�84z���:��ڷ̯�[����R����U�Uk+���ͫ��,`�g�"!/rF��.�u#���DYY^�?��ӱ�K�?k�� 4�D�=J�_���+�|Cy��{D9D�?��-���tQΗ���É�1������LQ�%z�K���OTWW_��tM�8�"��T��^{ۘ���ϥ�p�j���[D��y��@�_!HD=�B�ᯁ�)t��_C�V<��V{��dr�H�q���vλ<	~����epK�t0��INN/�Ȓ�{�7{d(b�}�]e��;��(�33��j�(�~2�����V�f�+rk�ާ7�'+2�����b�Ic��R..G��y�ngG"XKR75�p�ku�����&(��qSJW����ɚ�1M���Z�	���'X����{o��ߔm2�$��B��F������o_�A����x/���˟3�䥧Ӊ�>��r���@gBkΐ&���,�d~,&+xP<�5�ʹx�n������p�i܀�X�n���Yz�K')�(U0�����\�J����_�J=�Ʉ,їǕ�#�J"�N]j���L�����|����?Zdu�H*�U��{[8y`V�~
����a�y�Ƕ��(H;9�7�堣����YH�� .� ������S����ղi�W|O�8F���_l!���U�L ���b��i���b[_���Ͷtʻ�R������B%(�mn��I����c��ؚ�[,EZ����cf�>��SRRr�U�.�3q�'E>ί��=���U0��J}"��x�U\�?T�A�M��j׌����o7ye��q|�n�ئR�6��[[�|k�>���}��_�5�K�N�u�v���\V�'W)��5�x+�����^�L����:v~~�$�c�+����B�]�l�mN��}+u�wm"�n��b���qy�Gy!��o���Џ���Շ3p��8�@ɯ*P��q�@2,����f�-�݌u�� ���O���X�`]V��n��O�\��A��c�ҴV�1p��_�/G������xq��`҉��"'1J��r�~��D��C����B���)Uq!�


��?�X2����$z���^�o��"@���Z�/�>lhH"�Y��Y���x6"�y����v�W������'fi���g��m�<��S�8��7�̕�dv;/��c�����}�E6�'�@)�Uw=�;c�*�&��2����� 
��A;�nLʆ��`
�ϛh�������$TT�g�+'�*7�P�H�3����E�<0�#�'B"����=��sN4��fah�Og� ��/����c����:�;��綵�m(��梸wz����Mπ�Q��������������+rr"@��5����ɏ�b���e>����Nc����!	g�2m�:������"�J?�g�%�`�x!�A�÷821s-W��y���>Ƴ'��&�=]�:��f������'hb�l2x�FSs~x��$��V����&W:�֙$��~�E����#q��bv����x����Q>c��m69k�;?z�ld��,ž{~�L���C��)J/�v��a9]�Y��§*m�!u�z0TI$/����!����廁���"8�ը���;�$r�/�!�L��i�8҄�v�Z�!�XKk	�(���"y
l�4�����t��)J����X��P�"xo�iD��͸���h����djf����C9�.����3�}��c��j67�OJ �Z9�!	�H��,X��R������]0A�͙sjt}
K�b���L::\I�4$�*�ڒrwԛA�X�OX��z��Uâ���L9��Li^��Gg	��f�M������XŹ����CJ��ě	6Ĵ�	|:��;���� �c�oht1r����Gw�;��z�+�\�l��H$ܦ�ʬ$H6����<��Y�F�i�+{x������q�5��-�:��>M�J��	�'���Qw�"d�J_��&�����p*�6����u����W�{���)ծ�x9�-Q��U��m��o�k��#�\7]J2��hD�eD�����?��ֽ���C��X�������.���:�;l��}�dU2Ǉ[��oRA��;����\")��`��%4�B�;-�mΙw+Y��B��ze��\�p������H�c+�M���l�u"��Ȼ����w-���N�K��d�_�}k�Ά,!c��`�Q�V�KM�	g�]�.���~�^h��7V����n��z�馁f:�8���v���Z�Owr��{d{�J����Mƕ�G5�����6�s#�U����D�������8�k��8&�p�KWzcޔ�f/��\*[*.ʺԅF6U���ɛ�]�7���u�VD4
O��3���0v�]dh�g�|B׍D�c&�pv�M��đ�u��8@\A��Mb��S$Q��th��AJk���b�E�{�5�2�]����0DZ7�|������z���ߏ(�¶r�D�7��!0���F.���bs�8A��#ѯ��_��
�x��p&V��0�ND"QD���N#�ۏZ"�ʋL(ڷՏ9!V������$�@�q�<bһ�.�_�;R�l�$n���Է��qbuqq�`|z>��a/"��$�p{��#�1H���?��mp}��������v84 ��u5˚�OSiG]����_��eR��;��Y�X0oM��*�6>�U;�뷁��e��b��J���-�k�Zڶ Y,^y���ɫ�A��yL� ���_�߮��vbu;t��,�ݬN}Y������K���ak]�F����fj�A��Q��Nv?�ޓ���_(캗_��+��dmt��b����)>�~�$.r輫*��z]݉������)aˉ�X�)Z�ɣ�s�dc��E��5è�\��?QVģ<��-%�RsM��*^ybȸ9e��U�ü6W�c�D�w������<c���ڄ�$T��������s��C��!�� O�7�y�(m������ZX9k�>���v~�P<:�Vz�B��Z6�r�ȍ��~1". U�M�d19�l���\l7�KRn;�:�f����O'��9%:�&=�;[Y��vd��{n��~$®���x;	s���7q`��؉V��0Q�m�gu�^���?1�5h�ʢa�_��։�Ly�9;ǰ���!����i���^}h�pq2,m"�ɮ7���+������Epں�e�"܀��j{�PC���J>�oz�0X��]8������R�|J��n+r4��F��b>�qgk���k����Ã���@�|�Lx�PB
�wv�iQ�F&D�!p����L��t��U��i�U~h,'@���4��)�x�A�G��E������UV�{9җ��H�~����u�$@ko14�!jY_a�p��ZI*l!־�D��ؠ/f��� �Wg�V"���`�/��j�kz��`�a���
�G�s0p���'â�řR��o"�{��I��)�؇ u�_�Vt=c���?��2߂1��F�D�;&$C���䴻B���(�9�n&)�xs�#9�����?{Oh="_`9f��{"�=E򕇝)g	&������q�|[���{B�wo�/��2�Tžz���< �VF�$�5�.��a|�%e�q�,��Б�i�iB��Z6���5(YKV�����U�׹(À��,�xP+���Z	�q��g���d���T��T2��� �P��X�Tl�Qh�S��%l#�vZ
�u��h*�Jb��X��i~�T��)��G�����{��ϗ�Ϻ#�3�y��*V�ޮo>��T?�p�;��B�q�U�)Y*����9A�����	Ů(dL|��Sr�[���A�G�⛀��&�/���7:��	�*�34��G��*��L�d2���dɘ��p|���ld����Z��{��i�e,���C�2��@<"2T���/XA-_IB"]��k:	��,��)L�&��
�`�$FF2r60\ƄΓ��Kg�O"c_5D�� T��,�ʩu��*Б���E���h,蚜��yp�Xa
1�І�(^:l�f�J�0�L� b��"0�%L9o9 ]1��	��}�9���
tM]蚭�yBp�Ԡ���������[�	���*�Ua�:ѯ���F��D���7�-t�tm��C}`Cx�5�`��-j�E%��HǀjD�Hf�\آY�2��U�#��g�NK�CǦ�G��( f"Oؚ��#qÄv0!t���1��U
�֚*4D��/�*ĀY^U��Y�(��ǍT��b�B k5.\�'845��kvLv��W>����}���Մ�°Vl\NN���x�̆�!Z{�86�Pl,)�e9><��"�"h���p��#D�>��/���uR���Lv��?�Ċm�ɚ�,��JDφ�;���~+��=:>��_���N�*���?T*Ygr}?i��{�E��vme�:T�L��Ǝ/��a��U	��?������P��k��h�P�8T����Ăr>��b��p�T4N�"Ƥ�q~��7Xj%��Hx��%�퐙@�՚k������'vBK�R��6{\��I��q�H�lh�=xı��E4M�+䉛4�,yÝ�
n�#{��"�1��ό�9R)�\��X �j>��i�F0.��9�$J�S:�m��.��n�)�@�}�N�\�ԗV��J1��	)�N ����:K ���s�	]~��/�Jk7�t*�<�
!RBQܲ ��uvb �����;����OLF")�S�M��$��U�,=(�i�_�`�%W�+� �سy���Xٚ~{~�,�vI�<�=@�.⊆	��)���ЯLC�~qi��ǡ�C ����p�K��i���W�)��;���<��8['����C��%t��N-��zMm#��϶Q��MH��2��T<�α�И��Hs�}�	;8q9w�~����ާ<v�����QW�@(�N�w�<M�	Z@����!��l�_�@ri2x(��H�L��ڨ�$$[/��cg��	=��'| �͗����]���8�}�d���y���&>�!F�)�NN'Ԟ ��î��G�R�~�z֘"N:6���6>X�����v�:}
K��������*�D��Bʙƞ�^_��Cz�>�q~���䙄�^��>�ʵ�_Ez� ���z� �P?,2�{O�_혭������70���	7���ށͲ	ox(��;~�� �ꨥ�FQ$Ik��9�~�Җ����% ���;(�a=�Ҽ��0�ɍ�M�����u�[x��<f��])(~�rM*Ǹ�W�2M@��S�G���}P�L�o�+,w%�mu�^
�:c�4��ဏ�?tx�P�J0�v�_v�GD��;���7�x̎]�=�=�>H���[ͺJ�m��
Q��e`!�|�쌍W��H���F��B8�n�Ф�74+m�Y,�'}Z�70
$�6��O�C[�ͤ��r<���A����]�o�9��m��՘'����4�5$j�<�JE��c[J5�M9�oId~b Q���QE�֜]̈́�~-��o��\T]�6�1͕Z[q�b�$�"�=�rw�%"o��P�d]=�עr�~jv]7�i��3Ncr�ӡ&`?2��;�d����h��*W M��a�,Ǩ��om-� �m]��N�!� ;��=��£ܮP�h���� x�p��b�߁��j+��C��+�	�{nP�}(?�Wc��(�e�ɈEL��~��C����1����v��Sf��;u,x��Q?�/�]Q��r�GFPEQ��4R�	5"��	��-�?5TlP������#�G`A�|� 1��P?�w��&o�����@��4�&�5��w����d���K���7�]r��C��?n��w@y=mN'�`o�F��I2ॺv��d�ȁ�O-��\�!,`�GΆ
��v2�㈡�@KE��F���J(B[�\>cTi�R7PR�M��b�U1��bj
]..+�o���Ϸe�W�����z�?YA�Q��i۱��E.�\���1�����G5�+��f$��p�������m�b�����:'���~%%0�Gc��m'|���?W�BL��ʥ����9�v��;�l]���q޷������~�ތ?NO���V�Cى�|�{Z#�e�*{!g&`-u��SI�}M�[�����p	(��d:�wVds�C��%�s��QT;�>H�o������ �^�A���&%��{u5:�LD�)W��Q�K��i�1;���yV-w��&����|�j��J�%��fcM�A(�W/��A&!74��L���޿J�m��^�2�ͳhǢ�O~���{[�(��f�0�.k���ez������e�+�Q��
���Ϫ8���+Ø�G�MNn�Cdyo "�-o�b�ܰuI���u��"L	>s�pI��R6�6��!T-�r'��G�(��ZQ�%3	�vi�li�~|���/v����~I.�*<�r6X�+�s���,Y�v�cȘj%�7g�*"��CG�#��(����@����-�jq�X�ޛң���-���ȷ�.%6���n'P����я~�$�,yM�}�X@� z�s��k?�-C&{ �^QÚb����`wn�|�QN��o߉�u�$�T5�IY"�Q���Mc�}o�W[�`�?��ސm%����h�-�]��hdEt��~K�$��vx��+֎�w+�ް��4��tJ�+��Str���t�F�y�q���C#6rT�@�J�ş$��mΣ�6��>�L�S�D��Q@��9�U�$@�-�v�cJC,*u���fۧg3
�(��;�.Ń>��z���$�x�gW���[9Ky��1f��o�{���b~����;��%	��X=���Ka<N��D�.h��#���y�ļ����^�I���g�ׅ��*�@�_äg�I��`D��k'OZT	�@�t�rSaSX�;ė�<@���$g�"����C?~�5&��ڣ��V<%��e+��̳.��P#xY��F��(�_�˰�uBFi��j6B�?�6��'�?@
�����91���Q?(_��x^�S�I��:��b%_����;�6Xٲ_I�z�֢���~�w7�����r���~��5�K����}$*$��>�D�ǽ6z&7� ݙ���(e�~�b�M�)�����?��Xi��-��R����	�ݱ�5K5��*=�~��DdCV����1�9�a�f_�[
���4醗}΋d������h��,�Ơ5�"鍻'��X��������.�DG'R["�aҰ]���P�JF�^�Z�׆�З6��5�jrW`%�#h͒m2w6;��+0��<�	Ѵ�k��|�<9>��H#�hi�ٻ�@�{9e#���z��%T�����4K"��hn6���#���t�� ���ӓz!qPNy>z�'Ⴤ�VR�}6�!s����j,;�Xa�wZ2"eqH�R�SJ���Go�	}͉n�������))h{����k2���Ȱ��.{�'�峨��j����C�ى�r�o.G\��I�8��,�^���	I�o�?>e��ڹ_g�}3�ew�����p}=��i�w=�XJA}�iK���=!]�
��6TO����e��e���p_�yz��?���p��� l�m��N��|ο%���3��U�����Z�n3F/�Qy٫�.a��Uki=�+Ccp����	�*D���	T���R����	�I�F>[��OF�����:S� �#	IRj~��f�Hn���UAm�G�r֜�clT��Ɣ���7U$�sא�l���ܾ�r�Sk�$���� ���M;`�N����J���%�w!H��'}��(-��L �f�yG���}UTR��Y��r�h�������C]��V��)bA��
Ηy��Do��(�a5:�_牤Ə�|����L{�c�z���h B��Jv`�E��Õwv�(O8!��6��S�>���0�F��T�P%�w����>�TH���.��*_�����}�����fZ��Y몬۴i=��y�$�-����� e%%W�{/��Mw�N�������������$����6��K��"��%�U�TD[�M�~_�QIΫ�(,��m�冱����T*���ŵBq�A+�%ǑZ�g�sF�v��"������h�_�X@(���[�vj�|y���uH'}��E��{-�zv��]�q� �������_ח�4گ,�1�����@�{v��K���D ���/�Y����A������x�l�oF�����3lE1G"�t��C���%�/�k�Õ] Xכ�'p��?�忤����/|�yڃ.�8�lĨ6��).�#!�p)&-�`<�cS�&h��r�*�3m�ʵ������D��WD�1:��`����[[�̟=��-��Q�)�p�����Kbrq�!F��>�m��(>|?!%'��B��(��b����>7v$�B�3Yu�����Ž�ǘ��F�n�U�Q:Z�{��fM���6���W�y�0���u���{���ұ#�������{��w��B�Irj���Ht�Q,]�x��AE��9����?d̈́�h��s�@S$\i���P����C�g�Y���K��~�=;-y��u1��^�~{
�2D@���4{\�|��x��Nl���3�u�:Z������"M�h������̷Qև8V���C�ҥ�3�����N8�{�L��2�G���*p}#��S��|cmٕ�oS`O�1��Q��l�6�R��A,-�
�:��{����+'�!��~�3�4�W��/bf�*( ��Ջ���$��V��[O�i��Z<b�*B���r��6�᥆�+��7Û,I�cbb�oI��߈l� ����g��m'^FO���oty����ˍ5i�s��$7�3��JFX�l!�쪹&�A-��-�p_��:�y�d��hE/�V�f��VCx�����2����4	ȫKƸ�9aUD�U�mRi;|��Iji��}���o�XaoINq����'t�*�	!��I���	2��Y(��U�w�3^��=n��y���;�X�GW��i�?��֦�B��z�J�>��9@z�~�y�����׿���s��N%8TZpLhrS�n�7ם~��7w^�Jbnf+��f��f��˥5���"�qk���"md�(�VKeнф5/ԗ:?���G��M H�\׷�O{�B��o'6v�ǢCVZō1�#�.�O<l�8�9������
�'���wD�O�T����m�G������#�XD��m/���垆�Ӎ�����Ƞ�~d�	!�^��}>D��K����m�Qq�1�Į��K�6���AD�Y��}��'v�m�'˝�/SE��M�Hi��S���!���{'{�L��7��r/����r��7���׫����#�	��0s%jD�O'��1\)�Vfj��&��9� ?�o�/�wS�c����g&B_����&�;J�^������|
���G����ή�>XS����g.��2���|�GJH/�e��CJY#ğ3&y���Y�IzR�������1�ػ#���E-���a6#�,�拾�0zU�0�� 3���X~��s��O�2�I�� �!�O�|n@̢�����Ɂ��?�=�����r�p���+��H�U؂�-&��!l�.�j	�o��H��~cƟ1�'�i2�-T&d4�4ӷ�Ѥ�R���ƭ=��������]��E@X��2Fn�V���VІ������i�Vv\�x)n�ζ���g}`���p��{�bחʶ������HA�35~�E���dD�]��R�#� .��aa&���Ɠ$��!�c�h]*"��EJ�[Z���ׄ�lK�57�݊3�Ņ_�hDXPII���{U7>=�ou��/�+�LLVjӉhԬE>�����R��x��\>,Ҭݨ���A7�����E����8̛�Re��1��\~�W�U�\�a�
��^o�ri(p�_ř(jݜ��/~]4>��;�BS�z���(�I���W��S=Z'�r�kQd�uhE�l�M��j��>�Q�&|�_����l��,�s����"��v/8�no��I�E�W[�]�Mq�˄*0���v��v���eһ�}K!�we��Q�I3�E�1�W��%D���/5S<���k�o�H��#zi�(�Jʎ.��u�'�W�/@�6�jq!-93����������G��Gn��D̘�6rE*Wtj#5�`d�OE���P�/�� �����	U(��BRv���Ф<�+�e$	w}϶�IUGHSO�K �ʐo &�Fal�0��{��d1n���/}����C�#3j�3B�q�Y�"�YhP���4p��ګ5���D�c`�훏T��eچ&k�]礜��wa!���^���4�+E]kj_�M�.$�8�☊j��ybm��4e�e��o�����c_v/|5�)��M5����~�]A�����M��r���}�M�ܹ�eA�>���Y�MB�{��!�8����sh�˕u��2�<I�/%W��P�^�:d�#� s�H�,8����)@��g���r�q����c��
-�A8?�#��5(�O�U~4B��p�i/�-�C��焤;�5o7Y(.��eXc�1vޟ��x��Pa��'��4��%�y�0��Q�����bFkS{����i�2Ϫ+˦��Ĩp�g ��])�t[���!������H�)��� Ԁ�yI��N���ǒ�Ui���u8R�X�����n}���S�DŤ�L3�f5��wX8��_{~�G'�0�s)��|�% b(PoJW1Fj�_8��=�d���0�Iu���ݚ�H��)��Ϝ��wP,76�]�?n��N^,<"#Q�7�4����+�岅J,j��nl����U&����$�=a��\%%)>�'�d�KG�{S��$���ʌ*�$[M_W��[0f�T��WC�P'�!]g��mi"����[H�~7b�0�����5q���}C�7s=�Ֆ�ڟy�Dն��]#�"3�""��p�7��b%
G�l���RM�6���{���Y�O�=>��u�9�+�1�����aAQfJ��aJ�����_ ZEF�ד��.!��K���/��r��O����U.�NqI��6�;�t;�땻��%c�0��>̝�2�2<Cݨ�G1���јS��C�<5�E�(Ig���;f�JLW��[4�+����#=�p�j^tۊ3�� ��D����/��`	v�W����;�Ş��x0)��4/��B�\�.�4��_�&@�-�p	�ػd4���m��u�C���5Dz��tŔ?T��g�[J���Z����[*��ؾkM+.}���_���$��[̆m�|~�H�(�B��{Thvx/��IQ�r�~��[[��-q��n:�$�N�Q7���6�� i�3�#��fȜD�S<��Νy)�:�<&��M���s���zgtV�V�2������U3G��cJ}�������b�fiB.�w�����_5��O�`* �!D��j%�4��1$�3��0#ѝ������*os���e�;��a$��6AԊ�:��w�bB�W��zlj����0tF�4�J��(V~k��-��T�_�]�'�ͦ��G�-OfIeDT���\L��k[)�����^~��.g>L��Q�ةaˌ�g)M6����\%dnH�9В��e�I���G!��	��(� ���Ou�{���l_��Z�_�S!C@��u����:�Ϲ>�r�
��-���O*)��.�ֽIO�i�p�q�$��˾���,�XsZx�Г"L|E�������à��y7��'o*�5s�Sf�V/�Fy�9q�t3��?��	�%�?}	�=�����z �����������gR᫅��eq���͍|/VĠy�:�3/ �cz>P��_�p_v-�L����|��o����Y6,-��&j�8+ve��B�i��#q�@�i��]?{ �a�[���e~E �u�(RW9I�Wʤa.�Ĉ�:O1�li$��&��(a���J�����ٖ�	m\�$��<$@f	Οm[&�;b�换j����B�/���ET����z��pB�|Y��� ���X�l��k����'��[�H�ou�>�,�ON���'�8,[֐��Dg�V6D4h����V�1�\K��q��g'坮����W��'�|\����|X�	o���j6V0ii��Bk�������Mc:�z�%jKm���2U�tt�%����3��[up7~����(�Т!�QY3Z@�S<C���;��.�\�s+ծ"��[�)m�:V͛#|˕Z�ˈ�D�@>a���n<���੧jv���-���O6nS+�#ф�׽ ���?���g�0��,|�.nc0V�)�~(��t�P����vpk:)��tIԞ;��C���yK��$�bI�%�������)����5���-"���g����9�`���v1}��'Sڅ�`�ؽAW���� �z?�.����o�� Q2<y��
���$��'QI�ŒL��w/�7�^���GsD=
-��p��o�3��>W��J�#�^5�s��A(��@PȆ�P���F}�ˏ��l%��v#����a� ��R �$����}�2��ccn�=��82����^mu��p(�w)Z\�;��ww+���Nq����;��������Z7Y'�I�ܙ={�3�K)A}N���?1��h)D���x��Ev��a�0��X3lΟ=߀�[�����Â6Zr%Ybv|�=v."os;6ːs��8.B�3~b،cT��n�τL6�H#�e�[���'«q#�|�NkSA�XE6��zl%=���b!3h"\C��{6�'�z�In$Z�%����zt�;��t��o߽8��y��*��䞷*!�X�ٱ�*�Koż'�����b���)�P�
ee!=[�1�8��-����z{{C(�^����M����ި�~��\�br�j�t�sN�-I��`�����e��x��ȓ/����OT9�z@D?w��|9f�}���km��p���L�,-����	��Q���]�N({�*^�����Ći��9l���v�P���6�n��m��Mz	�N���H�镅���#�-GV����
ѻ��1	����[�0V�� ͷ�]<�y�0S5���ɂ���?��0Lo�ݿ���,'�#��v�Z�������[��Yb���<�%gZ:��H9�bl0{k���K����j�iS�+��E1v�����]�q����L/Z9����4(�}���!O]�|��o�}�'�� jgԆO7�)Xک�l��i�?*{��9�6x���
��E�Ĺi!�r�-��??�nsB�.7�&�M�D�Fl2P>�p8��j;�V�Y�.YBkJp��.E�]���	ҏ�Ԡ�G�hUqGk�\yt�s�-�>v0f	�B��֖��ꆸy�u�.�r�,
;��:�$�}>F.��@� �c2Tc��S��Ni)9A���H��z_o(�:= r�|P؛?λ�jLpi�t�y�^NT���n7�T���M�K�e���M-�>P��9+6�P�?g���K��g'C��ٺ�F���o�$>2;r"W��W�k��	��݈`���`�L�y	�P�j?��T�9v�k�֏-\<�"��ڨ=L3_���y���[�!��SG${�"�ɯJ����v�#^5]��5���&D�U<����i�r;V`�s�
��{G���
����0����ބ��L�g����|�2Q�v�����}��_�炃=l��>Gw@��X᏶�C�{�݋p#��m��;fy0�>יw�&O\Rj:=�0ȷ�u�~ϱ��3�4�̕+{�t9�i'��)d�v�P���V���*��ظ�̔T������D�eP��F#7�]�>���Ǎ�Dԡ�ғӁ͘�����'}��2�r�2LG����j����1i�V�?"ѫ ���g^+��{3S�x�M:�S�ܡ�c���n�Nݖuۏ�(*cy�+:9h��{�d:��Yh�@�Z�f�Ew�$�^L�tԜ]�XX0h]���SL`mOB��Cr*#�hbӏ�-�w۾���nQ^�f���J�{1>+8��T��ZZ� ��Xs��c�{f����X��7�9U�cC����Z��Z��4�URq��eS!]4Z�y�eC|��R��� `�%�Ƹl��^Qg�m9����T��	&<�&��[�o��`���DfL�;MK>��n���g������V�bv�y������P;S�]�jED�p�z�&7�_X�6P�1�;U"4�[&-G���Ӯ㺰scN��{�YV�Hj�FP�;�+76��kw~C�^�ɍ�V3��p^� ͕3�?����i�O-���Wh]F~��[�@�<��^�zG3?����Z0#Fn�ܮE��<EJ�V2�bs<Q.���rV��f3�"�L���h��1C��)�oo�{�3:A-��z|��JutR�cpd9��7T������]�ϫČp[�`�Z�_޴�;��x�wϯ�=�WV��r��L�1t�Rg��3��	xd����^�\�E�CH"K�z��=Ҋ�DHI�����d3>Xә�PѨμ�yf�_�16~#F=V��/P��0�Y��Rjؑ��d�ӳm���y��ˤ����O��C��O�O�c%�3�o��iz�k/r؈x��%���SY��v��̔=��K���o���O8j�FN���fi�Rᩂ!6x�R�us��\��l����w�\d�4����UT[׭3s~҇n�ŗ\|�?�E�,9w��/�C��h.�����A����e�fb���$F��֌_�Ɋ�|41�+%�����::o	�K�����jB��_&)j@m�e�v\���x��_�@������0�y���g �J�b�lٙ�Qb��e|�bTО5���J�H�g������0�x�w�D��<?m�N�yЉ��ӄ0l����F�����1��5���=�@u'a��(.�*�x�6���_)q��͛�J��j���[���4pbBZ�����G� ���d���f�v���dN��\}�("b����Dq�4�`��7C)2H��Pغ�����'ע�ƕm�\�c�;p�%*S���?�:އ���ο�ij�㘈�������Dӻ�����`�Av^U�����y�Q�3���"P�k9�^vG��@37���E � |ئ��v<J�e!�F\�W�2  ���	P���h�U�u\]�v,d� 9����j�3�|����6��/w݆GK�������R���3�#(|W�6l�]�#Dm�C����L.&��>�q*�?� 't�}VRB1v�oɓQrѻ��>cyz�.�v�^Ptu2�F����~�����h�G����~�����L�^M��F���F)��8�? ����ظ�災#,��A|<П(���PV1@Jf����? ��@���ʘ�?���%6��]��48�������0���$�I9��)����vﲇ<Nd�C@�0`6��$&��y�[FQ�f�����c%;���ֈ���@�Q��a�=2O�k����%��N��OҠ�~f��%`U����w�i�_����{+�j嬎������܊CC"��'62�\Lv
�iSF�U<4q,}�?��'��B�`�Զ�ZO�/'?�@���j����hh�v��rh2<���N�e�z0ꓒ�nTn��s��~��G�t(k4��)S�R]����t?q<���o#U�b1I}u���u2��87��8`��1���S����+�,zv��`SZ�5����2��c	��B/d`4
��퐷�/^�H�0
�7��[�k��,Ab�`&��C�с�i	�=}$��n^���d�~��B��������*�����^���	4P�fI�D��}B����"j�Q�,�1�5�"b3�,���Ql��/P\4D"7ȼ��OT�������uǄ���I:�-���X.4t��L�7�*�g�j�Cq��f`A���(���@����*]+�����D2�O� ��$�a�ָ�R��@�"��#P���b�d� ��I�:�ݮG��ɱ��\;�ܹ�\_/��V��x�6ٕ��1Y�x�?��g�֜%BtF,�g"u��_�8g��q�(j��u��Qjd��-u���6��Z�R�#Ip!��(jE�ǃE
S��p�E�m�vb�\E�!� E6L.�����`��_�4���d��E/�Q��.�,�H�4�n��!&�|Swsc�yV����֎��k�&t��hi1dT(<;$zL���j�ͧoa���]��Mg==�����~V�M�W��"/�m��
V9��1�	w���4��9EP��C���ÑaC������k���a���%b���Z�
����������,�!��EaJ�_+���7?Z�{�S,>�}�^a�k�80��ml����O#�b�⿏��p���JI���o�@H�YHrr�_[��J�	#�����$�=�޿�)���>���gP�tЂ)N�����͟����l�������Et���� bӵ�mp$T9��{��)U�X�ʮ�`��g;�L�VA�Ҫ�Z�!	�Ղr���V����`1:�p"!n�
O1�aYmu&��f|HW)	2�d67��V�]`�U�Q�A��ڊG3!! ,Z���V���G��Ǯ�'j�����m�ڑ/=9;/���V���R�瞯8\Wk�P���>\.1k��Ng��f��a_W�J𳮢�p��Б�	���`��/Ɍ�\�&X�L(fA���%�����WNc&H�tC���i��!2���Z��r�Z��Y��=�l��.�\�+��-��$ґ��6�_��������b�R�;ʾ�^'������*b�#~��9��`����g}���V���HF9.d�����4}��[mgqtt�Q��?�9��ɼ/(赵����j���.��ʌ_�mİrZI�4�>��;����<_���@E[n�ڶc�m�
ϳ�f`��p�F��~�3[]�=m��[�d�"1c�;�t��l�����c0���������^����/Om;%]LC�j,�)O�����z����Ԣ�#m+�<}n�]e�ބLr@��Pf?��l�U|�<��1����P7�}c)��O���C�5ttI�na	�.����Yr3et5i9�o����'=:Nb�����s�3���'0��^F�^D�J&�E�{��K�6���[�OV�\�������P�Hez!��*Q��'�\���P_k����ls�o/Pb��͎j9�E�S��w�Ck���=����٣�C �iy��f	`�pP�p4FJ����lU�������7�g�r��L?��2g���������p��*)��R�)fAV��8��Fm���ݍę�t�ޚ���!�'rc��8�y�k��Yw`o�[8LC�)N�[���� �.j�]h��)�\���'p?�`��A����B�%y$�����g�����cT3ɒ��*��d�Òk�ˍ�1U��xl^�b��"M�r�Z���z)S];�$���}|��1�%��GY�XE*TH�I�I�z��N�w��I,y<�6�c�j��W�b� �*�x!�C0ʦ<��$�f�3�������z�xVC!��rЈ��0����$�;��͛$�50�ǋ6u	6��"K�l�梍 Z��f�^hF���\�{�݇���J�
W$�p�Fܿ�j�3�9�O�v
<h��5;�^l6�jG=�#�đ����~F�R�]�
���?�͓�(��w�yL(NY��{H�b0l�2�!�!��
Ж�]YAr�ǒ��(vG�s����}'���/Ex}�r�HTU���q^�{��[�"c���'�?P��;f�/�SY�_�����лv�t`�j�4ج9����+U%�,vȀwrd��Z
�~���h�H�>e+�� 7�t�h$�.!73�}����ľ�"��q�xí#1]�������Y���u�������۴j�C�!�~�������屇���r!�9�7YV2��p�M�T��/�"��yն��8�Efn�>E���2�1n��� �9Z��?��v��U������?�Yv����Ax��G�x?��.�6g�21,�bi�e�N��B��T��:٬���R%F*���9˝՘�G�d'A��dH,���dS�c�)�N��N�Jݮ�����B��?���6S�6R1�"t#I*u�<�a;5�,=�h��Ѝ���
>!u�z�Hȣ�2T��ڊ�p����]�\�}��\*���jSܴ��� բ��Jv�54�(��ڔ3�Z{03���8��	�~���#���N��V_��r�ӂv�� (@=�������n�{�a�|�$��t"8c��3"Dָ�-{8*��u�<�/2�(B0d	z+�y��Cn11��9�G���uؤ�f�Mˊq󐺀���о��L>�#u~g�5��'����m���:4��G��m0Y��k�_�_���<O���j��ck:� �9�fΝ ����]�!���0�~�l��u��m�&�
'F		hT���?=l�J�O	4p1D5�g�^�M,��m����łK9(����G�*X�!r���Z�zަ�c3X� px�� M���������G6���t�~/�Ux�빗�D�õ_<��c���}��*�f���o�����V�!d�:k���#=��b���⬽d��}qwG�?��q���z�=7�\s���pa>���yic��2���}o��k]����<M���E^G�$���l$_hp�?�äa!�x������`�M�,hm�=�G?\�	���|3{��A���i�#�0î�����q��Q)R1��HG�	F�g�k�]�oÚkٳ!J�F|LF2��l�Y����f���K�)?��v��	M�1V�;��7��XhYo�mP=�i�۬=hXC���$`
�(���	��~.0e�2S1h������";�Q_-�	�4T��}��b�\[$R0��H)�.kB��V�j�3�jeU�b��T�ɍ;��Pg�4mC�"�_��x=o��:k�"D(ɶ,/���Zѕ8JY�4W��\���� �6�����y��v*�����L�
 �r�k�������?�:Q�mL��w�R���HH�\��K�]��1o5&%[����D���~&V�������h�f��΃�i�йSn˄��g����}�e6�Y���ˁ����l���k��0�q�d�ď�:ÿ�t<Xz`螏�i���U'K�~�����ss���R�Q0�,�8�d�FҦ�����gw�Z}��Ai�٢SkQy6`��̻�8�ٻ&E$ɱ�[�q�V�!��q�� 4\�f�v+�@]���_�*�;��b��&�3I�rw�^8%��r*{��it9�o��0�����-m[M���w;�?g�Kψ���6B��BUZ��bd�	H��yc�s��*�?�.�}.�_^bT!��
�2���:^��s�Bl�r�� ¢>�\f�]�k���,���Y�&E5r�"������1��b��b��P���z\=�ծ>鳸�X���Uh]��f� ��qxx�b D�i�%�elDA�[��!�����!��i�|¤e�s�4f��XD\<^:	چL�B7�bd��֦m(H��ܙ���n�v����������vi��o��Pa/b�'�zI�s�B'w~.���t�o�,)/M!>���pIUS�יnv/3O�S4x��$����	I�ts��g�;o99]�*����۩��uIOCH��m�o�8rW3��-/N��D�L�~7��������l|S�ũ
s��]�7L���! � k���� ֵ����ID I���g�Q9�P��˿7X�;`�;G�{���O3�L�_��џ5��%���P=�[�rq�;��l�<OĜ�t!�Ћf��ٲ�S=�|5��qcA�Z`�KXD:í�1F0>T%���4똯�6�8�7��P�2M�����.FT�y|�����`3A�]M��KpX6b�6tC���u�dH���;K��9��������(x���M�����B"x=��I�Pl�;p��\ �L~�X���^�KΘŭ�%]��1g=�緍4r��rjѝ���g��9����E�GZ햁���L�� Ka!��Z��p:��ߍb)��������DG8���fg:˦"�>7��k���r�P���K	8f��{8\�^S���f�W�,�x�K˭P���H	�@5��9[q�]��%"��E�'w�V�X�o��D[w�nҨ��h�ݹ�LdzC�����Oj��|;�X���A�c��Dm�e�[�|�j�$�TCE�4�� �c�&�f�L�@��i]^G�{�C
�뿸�W<_J�#�dK�g�5/g��/b�&���VP* yC��;�l�HA`��S@1=�ՆL�e�gc7��v>��`{N[�a����jX��M�{�+�2�8�dg���-Q���)_�����W�zb�e��,�����:�r^�5���;�
C�?��ϰ$���4eQ'K���c�_�*��K�	�G!
�����ô��P	g�S�j������
�A���5E��B��;�L�7fH>1��؍�%O����˰���zSPg���&���ET/���p��E#�u�N����Q�&&P�I��)�O1^����V|䳡�e��muq�Уq��R�0��ʰ��+��ҥ�)`�]Ğj�bO���f�6�N~�f�u�`��ui�w�A�����A��m�6�CH@R:O|��_�Kk(M�k�ά�zRv!��pd��~`�~Sj�'C���Mq��Yj|�<��	��5��9 �m^Q\�LbwvGm�}m"�,_V�`��~�9�����rA���P���Y!HqM�L�.��b�g�j�P�:��L���NsV���:�R�}�Ψ�fe~n_����X��̣�z2����@s���	��k�N+��y�����M*(Z���tN��m�?��y�~1fd0H�^���^�Ikm9��1�=���1��g]��%��j�-�SY���ę0��,{��1W�3�C��
|E��s`����9=��~5��&����T��)�����v�L�r8�MB
�U��#�~���."�.��2��4����G�><�A'��p�����DC+R6�$p� i�~).���Y�'K��H�'V��v: �>�����u��@pr�.�T����&�Ўg�nA�qs}���u�,2��q�1it
Պ�ȥ�2�/jcq��hy�$~��9���@�G�J���K�������e��a��	8J!s���n����H�4���q���N��֑Y���y ����W�z	��n�W�l�������L���|GFU��{(�:P�I�]I�+z���c9�^�;h����|k*fx���6��r�0��Qb���B�;s>��������t��C�lE�P����UIZʣ^����#G���C�g��e���:��vb��a&��7�o�"�G�,,c��;���T0OZ������G[���۸�x�}Ӡ��g'TCD#D8�����9�l��/7�+�,'൚�Cy�r}xpi|e+I�_���MC��v�X<3cH*�;XA^̎�j���gr��D����s��L�鄗��D���k���C��~�97�qbN�W?DĒS67��5�w� ��0�uy!4T�/��b���� ����'kw"ˮw�����g�KF�.�E:áԹ�|��R����y0�T�ώ��4{y܁��zk�8<��󚸑�;"�}�a��U7ΜDLmD�]֟� b6�"'�W�+i�t���:��V�w��V���f��q�S���׺�O�"��6��;���:go�,���V�+��t#��~*����?���\�<n*MkE�	�{�k��d����vޗ׫���˵���q�@�W~Hu��1��)�hrR��VV �:3�e���Z�j�lvŧ�s��#�%o���U��}���S����+�N���Kt�)�?z�0��?�M��v�j���_���y~$����o�߂�}W�~�Q���N强�� �cy!��u�"m6�:�ԟ������`�4*2mD��3+��lo�qa�f��~��(�[��/k{��|a�R��y�c��"�
�rCw밫��Rh�d-�Ѧ����ve�h���~sb�l6�/�#,foÓ���<x���36��+��V��l���ҦbY�*�Z�>�R��!~MC����g�ԙ�uC5;V5h���𨿛���4u�ӽĄxLC?��4����g���c�rn��5����ݬ�]�7Ý!.��(J���T�vD�#�8�2�ݢW�,W�H!�|X��]�x?I).��������m����ڞ����J\�@;�_cT_��C��F��k��T�Bi��_	��wMX?�h�9��݁0)@��{�<vj?k�!|�4�IM��!�hȏ$�tB'�u�+X;
�(ӽ�����]��ܷ;!�2�l���6B�MO�L�P�ʬ�}�V9��g��r~:�S��PN��z��9m$�L��u���W��"V�D�w�:�����T���
�Bk/�L�ґ�ty�=�D�rBa�'��N��Z�j����J�C�d�?jH֜e{8Rv/�'V�U�A
�O{F��e�;Ĕyx>>x@!��ʁ��|Q�hO�� $F䟓
��]�t���IE�f�:�F���hr*�,qʑ{)O~�9�#O"z	X��Z��*�`݋Ta7�z+�͗��g{��җ�؋��КV!-��ҁp's��|���������C%Ae��wA�=�Bo:�z�Ɲ�}��K���b��^T�4���ٻzں��w�P6V���\��]�ñx)���;<blȵ><��<I�J���5-9;F��BC��o��:��7�uD�ۃ��x�D�5[�}�O�8�͗�E:v���\����a��3H;�|�rwU����-����C��M�Q�tKa���XM"��I���1�Wk�$Cۗ;��v�w56H˛yjۇn�}s8�Ϗ0����v����fw��z�N�zh�� 	X��x�M����*�̓�+T���(\c9w4�u/���dˏ0�P��'��p໌-���Fo�"���J��ց�s�A�s��}� ��-{��� b?���|�m "�1�A�}���U[ ��@�J�s�t���@�����3�Ƣ�D�B���r�2��l�P�"����6�2�p�'(�� -�rYK��r�y�ԑ&��j*ܕ6�Wo�]��6�@�����"c����óEp���>ވ��_�����9�X�4?�äg�GAA졁��&��jQ?$��1�D����ו�9�]؇�WN�I0�{{,d�ؘ�/�x���V���ը��7w?`Q|�@�m<�p�,�nOX�%�s=��b�"�aY����B�KO\%q ��oqU>��+����d���X������Z�v�H`�-��):�3����,Z�Er�r�$);]Rn���4��3�������u�tF�uwJ+�i�q�mD�jܯ��_�����NQ��&.C��h����p���O��%����˵��U�E2���VOs������}���N�2d3�����A����/|�.��y����N|;�+�ȳ�Z��!R���/��E����JaN����x�fg&��cK����ܛ<��.��tƪ=ļ������S�M�b��Qs>X�|��T�`a�_��k���7�����1X�����{)�1����h0#���f#�����]>���L��Ͳ��(����^w���7Oy�~�Fd�i����x/-� 6�8e``R�#<��-{ܡC}j����E8�  QX�+% u4��徵��� Ş��Fy�ss���8��q�����^YO d�Ӂ6WQ�xP�.�]~A�v��N;.
��~�m�y�iک|�v�rE�L$�Uv8B.�� Jn*�c�g��V��<�	o���%כ��wOȏbh�ǹ�F.jc�ݻ���;V��g�;�������]�_�J����GF���c�g[H��D��M��";I:1]7Mu�L�s� $bFZv[�����+`��d(������;-�S�"��@�I�QƖG�#ʋ1J�`!�T��Ґ�˒�-�˓@u���$��L���7�E��iU�f������*=�e޽_���Ȼ�\��@!���I6b�2���f5�8G�� 'I�p�1i��C�%Ռ��s�������v"��,և�D?�D�R��;��a�$��@��� 8�/���T�c'9w
����p1K(��j�ʅC�"�M�j��o��i����s���m%A���1�Q)��9��$���L]��dX��3)�������4t�BO?���[M��я�����S��m�;c��!-�MH\S�&��`�φ1���7���jh�o���Y�˹����G��<����^W$�AQ������S-zF���.�w�ԖG�a������,Lc�4��S2��gF3��WyT��J9��;���&T�6���� �c�`��;�03��k�����ړ��*��a�7�s�Į�|�wc��J�t}������ʈL�x5z1�_I�v�������SI�1+�o9�Jb�;*�l��T�9j�Z\wr�$9��v��u&��գ�t9�K	�;�; �c��`.�H���:L|� ��`:�Z��<���7hhRc��\�5�^�
���(Y����X�d ��>�����(|U�RD���ɬ\��)�ޗ���z�b��X��1C�p�B��x��ĭk(��<�����<63$��_��D2zTy
J]�[��^�)���ZUؖM�x1���#=�H	J��9�XD6���f͓!�s�m�#����a�G)�����14����o2��-{�i�acVc��}��	��X��Ea�a
��&�XNR=#S�o�[>�*��amxg��//���^>8D��~5µ.G��1u���t�����j�hj��#���M�X�[꛱HFnn0g���P�:�a��0��7z���X!݁-?��%���'ȷ�|,p�+��lhz��8�+̥���oP7�=[���+_F�2����8l��l4�Ud�ٓ��~�-�1������aq4oq�!oEm���_���I�(�/1��⨛�0�	�G�7���Dv4N��YL(�v�9��4!_�� ������`y4�/%c���r͇hR
��pDT찪)��k�e����4���>M�#��`v���0fh�Z�&��l�)�0��qp2A��X�#��u�k:/��Ze�Sa�9��;�m��������~�>�杋����p�$(HsX=Ey�����%�@C�
b���̖_[�B[7����'>(}0J�t���l���0̄�"�й�6D䩔m�F�j4Β��HvuZ������I+�4�7�^]��A�'##5�7O�M�T]_�d3��6����#8�h�Lou�NE(O��Ɨ�0M���3W�S�,��C#=C}5�ȇg�8��R��9�rC?���KE�V���2����w.�>3�g���#�X�E~jnJ��r�|��.e����b��n��_4�<Y%��۵���\a:�e����؎��_�M�Ϟ#��o,���G�z�(�� r���	��
������?���
,���@VZX~[����T��=�;�kl5^A����.�0����vR���z��:���,�Hx����']̜�oyK/e6�	Ke(�:҃#�i�ҲZr&�d52Y�7%����[ǽ�N��_�-H���!OH�����x����C=4
^�\��UN��q\Q�9�9�iJqG
�M�_s�=�>�^���_�z(n���d=\�0���1�Q8�쀢�f�A(�aLU��,L���<H��ۖ@�+��P��J��� >��BAr�VhL���Q$BCk��c���XD���yA}�î���oݥ����i 1	�����`p��/W�LH�a�vϟ`�}UoS�4N�-�å�>���W�ݴ���H�B�=���"�Zr��G���y�&+��q����m�GylG=����%J,����fG�v����>�&O�_X�D̈́�eS��8]/���0�tSk4u^-`���&	�\G��Fہ:�b򨡘@�>8P����g��"4'��U4Q�AO�CR1���>I�|�_T�w����Km�*3��GI6�0\՗�Un�����ٔhՎi���y|?]ws�6K�|���k?.]�g��0rع	���'����z��osq��bl!��������_P��K�r���s�x�N�o�r�݂I��N�<l��S.�fΣ�܅�S�knWI��op���&�A��{ԁo����s��#=;%�:���C�<��6�h�b+}�Jz���
Kо�Z�V`��10���>�w����
;���$�s+�:����i|G&�W��V��D��}?-;!FW0m�|SC���Y|�Y�n���8"���f7��/'�^� ���ص�P�mnME�}P��XWK����\�ʄ�oj(EUc����m83��m��ah�m�������@�`(K��L�L���x{��e{�b�ך(|�p�N���͈ɧ�B��~ȴ7���oS�s��{œ�̳�$YO]5��Ŗ-�[�Z�q�d��;���(�}���|^�@��q�A���@w6�9����#Ux@� ������������g����Y۲�̸���:c�UM��²yy����(�~հ�����e�^����
���èp�KLqk�n��j��w+�1������c��˅v�S�Skm�B�)�Ђ�#qf��i�55�ѵ�����&Y���U&�z|�7g�4��H�#�!}}<.S��v�h]��Hǖ���Wb]]� ��p��I�g�F�n�Gž\�oT�!�+�g��܍"_�%����2��țF�_,�1Gr�<�}��xk�X�K���~�r(�d�	�{Y�ho��G|fN���Z)�Ǧ�#de9�\��	;>���f`S����EL��U?�S��B�7��e��p��~w������SU,C�_�]v���jw�!��D���m�9X��i�@H�WH��~�����m|ʍd�~s�#������כN��><"/ �m�'��D�$���\� �?G��̙es5;�b�~3���|}���Q�l~'o��|�����08*)�Y�%��@�߷9��{ŉ�%V��ƴ��4����i%��;�y�N/���:�8.^����Q���f8�� 4d9���I����.{��5����
\v�y�������,M@�=]��f���hy�ԦպF5�����;����uH����I���:bQQ�9N�����ß��|�Zo����հ��k��וu>���ǟ�h%d]ٌ��5��v�	�u�i`�oU���|8�,���v��|ђ��\�4�LUA ��1z�r���!�g�Q�I�6��I<]�����[�.�9ʪ[�����M�f�yÕ��q"�Q(2�F�	�����˻2���·���+��bv�|���X�o��a&����x��k,g��d,#�K21��A,���w�Y�J�l�PP������JHj��-f�q���0?�6i�'Q0���
�%e���Y��f�~��w�c���;�!e��3@l$�r��׊H�ټ;�x8��(��6����Q���Z�Sl��X���ؑ���;�����!��Tj��]c[���4�+�ޒ��d��b�Kz^�ļ�=^�#���qh��n�Cm��c�r�E3�<s^�9&^	R���UKo(�1�D	�����z�b�dI�$��j�����>��E��@�"�4س��r�X��5˺�N���3��b�����n�v�1#c�^x����r��
�T�����OP_>^Y���T?M�EAt��{F���֧(�~�+�� ��Lp�V�!
)�t��/[Yo������(G��8O�1��Vd�1���	4��! ��w�tz�t��cqB��5�aZ*�jU drBi8JZ*<�f�QԮ���;{0zSQ�1q_�%S6��ׂ!'����ȥ�P�q��۾֡���?E�i_��x�Y3����e��u�_.�>�(B��D�&�X�Aj/��$������TTĊ�|�EM�W����/	��,%�'Y�T��?�i%�P�}C-�y�8��[ֵNW�+d����٤�#Y,ꑭ>���2Fd2c��YݟF|����L:*.��b ��3 ��i!��S0�!��'y�Y�*!�ɑ$Pk����,�]��������|�T���? J��NH��E�5��E��.�>��Ɓ����l�a��Oh�a ��ȕ]�ќ��>M� J#}dÁ�T�00XE&@'��L�V�X ��P������X���d��:�O$�4��&�0@|����r����x'u�ǿc�dM�yZ6�z���fZ1�CI@�R��=I-T#*�$3>��
�9(a!��	uZr	�ʨ˱Fd!� <=DQL���c��>/�Ke<�)�X��-�_9�Mit�a�PkSjjLh�)r�K�uW��
F��R�[��9�G�ɝ_ğp�)(����\������Nw"�����Qfrg��7d�y��:�S�nt�� �=�V�<]���b��x��2�-�)��Zp^��J)�D��<�8UT����H�+�p�"JC>�Uy���A�,���b��PX�f�D���:�h��ݎ%�S���eG��jUQ�5KŎ�KV� ��gv3�K>T1E4g��ZF�磙~gME��h�$&n",����֤�7��ݙ����3�yz?��'���g�)�X ���r��ꆪ���*.���琐L5��kƪ-��:l�b/%�l���#Ʒ�P�N�[�*ʏ��@��Z���h�-�x�)7� �"2����V�L��/P�~+7���a����i��Ԇ@�����4��JE��N�.��g�|r^��g��î[i��'J�s�<�p�~��*2O�F���~aΜ�g�Θt��@����jrs��j���F����8�,"� �?���-�&p�"444 `�B���\W�]�dB�=L����*È˔Ýd��!	G���)�����G�;8G��[�Nl�۞L�L<�m��$۶mۚض1�3�w��'�ԩT��;��׷����^)z�d7�Zt�M��K�7$8���\B��������WF�%N�DS� �W��gˉG��k�fz׷�#"��dz�d�`X�������wM�ݑ8C���v�6R��-�=Z�w�jڻC˄��!q��@҅2����5�a,e��f	���G�z�oˍ@��"�����#���Ju�A}�9>..�ޞ��'Z8A�Z��tx���G��<��d:[�/u+�nԉ=����Jiee�d�8x���_��$�P���0�mb�!y�9A!�/�S�t�
���
�^$M�r�a��00 B|�k177���H
�%nh*L�v���T��dtl����RmtrS!@X�б!�;" ȑ�bM�(.-M�׸'	��K�L�K}�Av0�$��G"'���UW���LA%��eg�{�`G��-�����u��BW������?�Ч�4xRcLW��w�[|cD����B��y�� ���a �T���D�A11�_�Ӑ`� BHJ&����,T�S����НVſGW�2����s�ϯ�0��:`�)��j���)��Z�Nz0(L0��7�熌."4���p?&�>�,���O�x@���O�C����as)I��7��Ȟ��`�K�qN],VM�!���N���DC۪ʈ��$(H{OJ|�+fۦ���o�����5����q�˙���W[wnM��It�Mny�r�U���AVS�"(�<+�ᜃ�t<�����]�xu��������锭���s�p�"nw�D@�nS��SL���i P�3��M%:p�\7TAE;��jR#���CRwx?-dp���Zz̏&0�4t��o�r6���}<O�j��
���7������}j�NM����'b �YDpz��eӝ�����#��I+���;Pv�'�e��󖢥�~���Dڵ��41M!+Ɋ�?���5�i>����J�@�1n�������s7�|A��O�A� �O�P�-�k]%r_�ȿ�}@�<��k�p�>����rk&�ҹ��ܸ=:愶y��9�QL�-�,���s�(a�J�#뽆2ಀS(?႔��9�"Y�h!5���$��E����h�y��6���H$�(P���s�2��y���Xn���c:�y&F}�)kJ+�r����-})۾�O�,��2I�JbP�\]��(j'�pJ�̂������e�P���w΁���,rU׭�rx���M�,��AO��$�
�X����A������z�;���8c�g��-w6�(��f2�+��עc�3ݞ<;2�J��c�����)�K�ժ^�S����|m4�y��	�������/jZ�%A�bnU��	nJ����Rڽ׺����ng�O��/-���o�N�]	�'���Jܓ�^M"MD���	�ь[E�I���<v`�o��f3ny�9���3/���Sc�BfM���1N���4����ު͇��{��5<=�5ng�;0��{��/ 8O��v���?r���r}�����AwȦ �)�����`���=�ʛ���'̝1��J;�������:yH�ߙ��r�s���,��؛��ճ�$�σ  ��'�_D��G��@TQ'\�ϊj5�V�8����?��e$R�7^2n񻽵�U����[3RK[cI������կ�<�.��������5�7g*{ktj*?��h6��S�#_���9�� ˡ��;��D��~�"��JW�G�����KR�Q�z��+E:[d��E������,��)��tٰ��ӏΆ�d�~�8Tf)��uxh��I�k�q��4֩?N�c6��^\Y�u��]$)���K@5d)m�X�C+#4�R��[`�T�����0���H��g�S�!����r�ѶORc�U�ժfG�RLm�����uآy��T���BqdP� 4b	Ԧ_1A�:��$9�燀��L�y�;o��[o�Ȱ_��r�a�^9	���NKq�&�0��$��NmT�����5=�����M��y��X���r�saJ�
k5yM%���d!��5���`�8Z�.3��ǄS���H�P��c1��݌H ��nM���0�ڽ_.����[��W VȞ5�?ʜ���/�#zp��"Ew��&�cE���'�PI��4����?6�n��
��a	�"Ǹ(���="���H�{-�C���B����)�YO�j�-��7$�B#�(Q,8HF8�D�F8�`��R��	υ� �#3���:�q5�$�j�ҽ��a��tx�n��{�<^���QJ�@kw�'X����p@�P�3=2Q�O(Ø�0$p����������Z.�6M;��k��o���#; ä�C�^�ls;K%d����x��l�y�-�Fu�
�寴-�T/k{G�U��«̅n�z��-��m���L&!�Hǭ!'(U��)bte�#��H`�g�	ոi�����N/��(H��grњ�A��X��"�B�� ry=j�I�互�}ۢ�?@k��u	QBw�[i�z�;?UDA��N��N�l�{~�9�k������:>Z�6��I��
���`p,��N�ǻ�+����rWv�1��O��(�������3Ո_�u�I0+M��~�+B������~�R�y=� a5<*t<��D#*�S���N�;�4^�����D���&'�3��rN'�B�m�@�v-��rPz���0�(r(w�Ǿ�E*��W���3&~�Ab�[i��V���ѿd�m��a�b�I�a�J�.�Pi�^������m� ��s�t6WC:�3�!�m^G��lx���.�J�[WO���0�ѥT`(�d�#�q�q|���R�� ﻞӾ�{B��z��f�q�yY�M'6'�«~!7�&��ϔ�tCȒm���k�E��ԕ��#�0Ps�W���bbx>�V=��=�n=����&Uz}���5�=tc壼�wC~}��Q�ߤ~7���>�4ːW�7W ��E� *������q6��)A��A*���]�RV��~�JA�C'�9ߞ���rșW��U;��*T�cԀ�b���Gĝǐ�����:�fWo�N�HK-y���MMd�q*�忞>���1����w�pq�[%̞���#�_�����2ZX�>\
�w�J�3O�����)F�ۡ�UT3���<��Rf����"p��RT�0�+Lǭ�3����od�P�i��Jwp��"ֻ�@��N79�ņ,e����~��)J������v�xY:�&�-AFP|��F0gR4��$�ȓP��?YL鸪��h��8���e-��7�h씵\&�j�:k�*>��l�T����C\���B#�F�!6ϩ0Jh>N3��6� �H��nO[��6Cڶ8�F�JL[>���;ο�h+�0D�g��`�����@^�3�͞s��**���_�h��=ϡ ��4M}�� �s���a��LE���DNZy/�A��+~t^*f�ʇ4��T��.�OˎY�������,��(�E�g[C���4i�hl.�M����5O�����I��8��PJEwx=�gz�k�@�UF}T��Y�Ш(�� ��r�U�bJ//~:M�^�*Uؓ>���r��FZD�}K����9wmT2RnK�Ȝǯ� �_�l����ƣ���/2.��!����
y�2�V\�m�	[�'{�� �v�*Zl�?�����oq�K�|S)YY�ۣ뛛�Ώg��؉"N�)\5�)���b��]��~�{��?6��\RbC����
2ѯܰr�������ch�U�b�+u��8>�ө�� ��e��y�7�k%���s���)
&�@gp�ٮf~ُ��׍��xf?�<���.$���O\���b���ܑ�����)����{�T���yhS���yݢ��[O�S�5"�<y����딁ɜ�.#��Va����֪��
f�`}\���#���	L_�hEhŵOZ:T�7n�'�F�]��S��ElO�B. ��JO8����8Ӻ��z�a�����Ew̓v��ِ��*�z���~Ҥ�޲!Ve(����q����.=2&���\�E)C��j~A�Wւ_u����N��g�W:|	Gr���%\�j�x��s>s��`H�����<Ʈ�6�X��Kz.�	.S���&��KwҪ��kk��<��u�t�����HLy�����YN��]�d�+qԅ�-�G)Ygۓ����q�X[����G4�Ap1���w��B��O$f�9�-6Z��Q����S���1GV!>�!~w�POĦ�����������+�|mp�f��/�@��)�*�'�����$����Ĉj5�ua�q��/�,�Y�����\l��:�/ PU�j��E|c�bHK������&����㙞��T�D�j�)*��Z��^���gO#�t�7A؛:
�|��F|Ԁ�Ä��C��@)F�n>�ڄ����>����t!��Qw����TԖug�����X����A\�I"�w�tx��D��]V���
�4�1߲��7��h�5kt�o1�@��i��^�����K�\�u9qq�;}eFզ���*�b�6ł�I�i̢(�Cre�`H���pjۜ �@��qe��Q�`i^3�!�V$wS���V���{U�y�� �Zv�<�Y��"h& ض��\��|�{}ɼ3�%���avP���P3H0�Sj�A:�Y�Ȗ�{;ׄ�gO-tO��Nv �ݡ{����_� LϏ-\��XGX�N�"}��t��t�
j�X#�!7�a��o�5J�+���]�۰��:!{}��ۿ��k��vٷZ�-�����>��y��y��w|-�b&.Ī�8�٨�"	�H����b �l$,�G�
>��7ՍF��m���Ȱm�h�_]�_��Pud8h@�~��~T�7�e]�dltHQi��2Z� a�lU�1�<UV9Ȁ�^^�c��wB}/��,�~D�.�$�Za7sR^��uםJ'�cӾ��5`@�:��[�����[�6�x�����|P�& �[W8A=�e�	zz�jX�*~��HJ�
�ozȱQG	�G�X�Q����H��}#�ဖx�ʸ��Z�P�u"
,z\���y�>����mx��\��o6����z4#��ޓ�*a4M�s�xr#���Ø�{yu�"���CL�(��˫��LE�We���ؖ����39�֖�3u�s�YWo��g�j8���P?���׶|�M��c-9���Q��f��e>�?-�#����93�}LNJ���4tT"�����%��x;��M���;lh%t��%b��s���\���=���;2��Î�ﰣ��=�(�	��7���Ǫ�!:���Qs���YY�Es)W�毷���k�
D0��� N�����hk�ʇc��ks�>�� �Xy����`����]�؈�KƗ	����Z����==.�h��`�H M۫h3NK&�O�hOP�X�T�ގ����jM�׍U8_� zA,8Z8˷���}�RA��c���,�s�}�oi���W��-��e|��d�cmפ��]X�i�w
�.�M������e���I�:r�=nx0�w��[���aA"�|_2���v���;Q��O1 MЈYp�?��zA�"T�/�Dbx0��F$**�"V#�D�=LI�I�3N�XC	��@D	yE&�����#�πC��[iy��L;QG��)a��F �v՗�(@�XV�0JI�)�uM ��FB� �E������lЪ����`X�ӗPJ�D[?(o�;:�3L�7���9�O�0
�]C�1���Ֆ=}�	��ӫ��^��R�{��L�t�؂�)�E��k�iH� Y�Ux�
F3$j��u9@Rk2���ޓ��G�%���,)�Ë�S����,���Kie�8��v��Ap�)X���f��d�0��@����N>	�<]?�``��B�ŉᴣ��ܓ{�2K^��m������q��謝B�����L܈�ⶆa�P��߁xo�n^��6��<^���K|���}�݁W?���3�:�TH"8߆h�J�Wy�Tw��[\�?�e��@�w�%]�Tdq��'�QG��i*��ǔ��A�8�QDR���C�n�n�@Cdy�vݸ�%$$�g�\�ʛ�P���<=3�	D<(e���/9���<�(V��}�D2����L��rL���������(��S��2�GX��p2�b�셇�E7�/r��c�Y�f��GI��!L[��o�k�)r��z>�:�/4Y�wuc1��mp(4g�"��W��r.�P��/�M�l�2D��ֿ��EE~�A�+Lc���7��4{��[j����U��84���17�������y���l�l+ڟ`�����
����)"��,���O'��ε�PRo�]��@/W���թ�����?�vq�����sf2�琣�ۄ�v ��@����,�~Y{)���)��C����g6�J�qY�	P�Ы���r����lo�2�ϛ��,Qt�tA{�6����`���彤|@���|��ha���!�AK��h:x��$��$�!q�G����U˙��Մ��2�	�3��f3�K�z`�#;P���dmփ��qڗ�f�����aQ]���c�:���S�k]^�졟��M��P����D�[�B
��b��VY?����a..��-���ׇl�A?�A����0l�A<��2�t�6�}v���3-M�-O�H���.H�ޏ��ʫ��L�'�`B����	�$H�/k�|�k��`�XdJ�VKgL׍
85�����"�Qp����n!zkVV
��j��PО��k/��غ�ۺ�oۺ�2��1&벦������AA�� #<�\�
�b���!� �Q^��yP�f�g�_� �lE6����5�N" �3�o`�E˯"�/§s[?�8�)O��2Dã;ER�Y���R�'��Ƕ��N�R4����Eט8�1�k�3T�'����=���ꀈ���ZZb�kRAX�V���~%���$Mml����`l^lDA��Ht��!���	��͎�0��a�_����+���L=�-m�*��pÙwE�������0>v"����-�U=� ���j�5�ga!�s��)�($�u�z�i��0�����ˡ>=�*}k,��:0��V��d�H?,ʳ�MZ��� ��Y�pUm��:27+V{��w�����.����@/��~�Z�@%�Aѻ KRc�cW�w�ͬh�:�l�Ze(���+x�E�<�&M�8Ɔ���gp�7��y���� �ث���i���3�?׀Wؚ^q�9<y�<M���,�k?���te�7i(�AԲ퀛D){fs�_!��t�+��W���g5��
�=� ocQ!��N�~E�8my:k�Q<>�8������^]�[U��HI��v�ޣ=!c��	k�*-��^���<�:-�KDhg��G�L�|X��R�YB�x��2�#1�L.��E�Oa:�]� B*ߪ���]���h1���U�S� �t�5�`©�:���mEl ��ɫ00{�J�Ʀ��8�)G½k�(y�?����lgr٢�j ��w6;��{�4�L����!iŦ�h��EB@e��x�粷�c�5����5�xY�ph���~�awN�Vy���F���6�H#s�)�!-��(�cւ�O&�eۃ�e�B󭨉�4n#%UUO��`��E�ā�3�u@ �1��p4�U��^S�!ihp���r��;������cҼ���/{v��$]�:�H5��p������Zt�&$힤u�φ�`k�����%��+g��)��v�-R^P�*�����K���;�g�F���<��h�v���[���f�|P�M$�Q����|��@(�0����6�m�>���{�q7��И8Q�Y
.�o���R ��h�Bĵ���st��|�Qb��?��ߘ�{�.hX�=�����(.���::��k�s����[�fE1z���^>�v9=��RQ��/���8g�|��t
���b��@�x�n�����9w�]LY��^�5�iw���*��,���m���q-�RVȖN�W
��3��C�<�/`f\�-C)��qwy�B��Seg��)��q&��Pd���3�S�Em^˚Z��a��8ˌT+z�ĵ�
�h�웠�fod�}�e%�MC��zXմ�����3���֢v#�x^��D�L'�ܼL�-M�n��e{��`he�d���W��'}�����)���V�廤�p-�cy�AZ�*�@�ig���r��y���ǟx�2p���zjq{�/B_�`^�G��!�����AF��a�+�VM����lbx{KRl;���K1+��.�8��6L2��o))ю!���z���Ao>;��\L�X.v�nF=`��"a��X�E���������]xї[ލ8��_sB�K�������Y��̵��U}����D�ƞq0oU���T*�,T��h���,K�z��0�Fw�x��򸾑�qލ2�G�G#��Z�u�r��M�Q�"ybuT[D���x}��5)��I��,vt`�s����'�}��H!�~�&�AƔ���,a`�r��k�1��O��4��.����i�E"]<`������ke�#�X����iZ�����ܠC�\�=j�g��g��.���{�JO�c%��~��%`hԾ7aL���ep�����y7(�
��`'�m�`g��=YF҃Z4(C!�+�g�����/���NC_�d�Y�X<q0��ԵY{����%�h�H�qɿ�K��d7������ś�x>�_p����6�%�qy��=��RQ���Л0�|%�������ƛ�}�/�-;�	E��P}���3ѕ�������u],�>���?GV��_�?�Q���B����n�\�z�%�Z{Z�=��v��^���;���"�W=�&p�\csR'Uy�װy��y[�<7�=tJ#�t���ɍ8��Yq�K�D�(:7�~g��JD��fپ'�,V��|qdG{���[y;Vc��Ʃ��}����U@�76=ӟ�g�#V!�dw�y�����D��kI`le8�u!a����������GZ��R��-��N�՛���"u3<3{�<��QT�Ѭ�.��0
��I^�K%����K+�I��O��� a}��U�1�-�G��E�l1'AW�ʪD8�<�όe�Z��i��,k%��5��=�&���cCќ3���Y�m����ug1�Kw�ԓ\n����#����m�ࡧߔ�A�� fo?	�o�`��>�-ZHru��D��ޫ��J]o�B�T�80|N5�?�	�7��Ej��|�-����&X�a�>�>��ML�@8�,���]�I��ke��K�ȡ�����Au5�4�U1}�Z�z�#;zpB;� ���0�����Kt35�l�����^͚��D�>w�
���3���v͹NсQ	��wF�P#�w)	�?=���o�%x��z����:oYh��6�֛�c
qE5��U�`���2��y��`s��}�E9�~' ]oo�
�֒o��/O����RrʛI|�tXRBҁ���Å	�vhx~L)��[���߾�G:{,�]�.$_�$5xk꜏�q�N���*b�3��I�O�j����R~W��N�E_����@��c�^�ZFϲmS:��5�*�2|.��W�@pL͂q�H�_ݞ�X�"՚����g�1��Yį��F�����ґ⤎X"�;ԗB9Nq��T:��ј�5�r6�J� ��mW�VΝ��V_~���a1� j�
�� Ӟ�G���D��d���<L��'��F^�K	�;s�a�%�  %�vc;�{y
A��a�,�-�K�tZ~bQ�H�"s]yu�Ԫ筂&7��ɻ
ѽ����"�/�f&P:T����]�I-�.��y�P"���t���B\n���#0Y�F3��Ct�϶�AD�{dM���"h&��48�Q�q��s�,b �3OOI_�NK�m�·T����z����mw�2c���	�;�%���s�9�Z $4�+Xg��D94�9�RM4(�Л_��?��3U~�x���J�밅����eb�4�dʀ����;�	�yD����U��(#7��[�(��f؛���
N���9�ԁz�?k��Eބ0U��]H12\�⣔��vf��X���K)�.:͏�7�ka_ӊ#>'G�a�Iǭ`�|n0y;oH��j��"��㎯��v,a���]��N�mc�}� �#W�.���
P���S*��ùD��ũ����rdQx�^�_)s�@��9��:�?�*y9���,�Y'囡��ņL+�ni��k?���O0��9�y�?�^�@q�b&9��4z|ϻ�GW|X����h�^_��7���r�k. �TJ����ke�af�y�̊���ti�,&1���<��Ac�����5��v��o�N�v�WkQ���u�m����*-�ɬUD�˝��`��款C����Q���[.�������rh�Lt�-��w�� 9��dTR�!��%A+�Cڗ]Vْ�B$�fށ��M��)�V+�ua���{��5>N#�Bqee�&��ZH��~Źa�П@��[���
�3�.��xe��;����wwo��)D����8B���{Z��N?:3�h�x3��pn�rC{�TZ
��Fy̍��RD�ϱ�6^�����
hX���P_�,V؝��'���Ʀ�����j$�3;�q���]bȊy]d�\Y��+���n��hq������-�E��c�Bͧd��飼�H�Ƅ&zo�� To��"�g�L,��X�)�Բ
h�gn`H�y��<����GR@։0���+�"î"��P��I
�X��܋�=��0����9%z���y�m���k5Н?�23RG�V`�9,�?�L2/U\����49`f+��ׂ[����tQm��:�J1�9⵪o�S��߲�:���b�AT���ɟ�%w;94�K�"�?EM��q�����4�����6tmx�Mt������2= `�� P�jX^ڈZ* 3k���TDd 5Ԯ��t�S��'v	�ei�|���������VNQ�n@�n���^��=���զ�Ǎ5o��ea�&G��!s���J|����{��)�F�8 (��,�/�?eWhl��ZE8/�v����I�r�}%]o>#((\�*#˪V&{\z��T���%N��Ö���ڱXp� kW|jI�\�0T!���R]���t3`��		C�y�����K�2�A���%7�[��	��ӫ6���;�&Ƴ�& �="(PZ+���\�-���5;nZl�#� ���ٯ2�:��A\9`��5�<�Rjꬻ'�Z+�o�������S>~�K�Pkפ�K���/���q���tހXk� +t�����BSE%�r�[�嵺�S��\��C|�K<�Q��E6�lGT���4N@�SJF.�?�5��<��|j�W#Б��sd�x��r7�)�To	�h��+�'U����ipf�oң:@k.�<��[���F�˙'g��J��{ ��a�\8)/��j�l���-��Kd44�]�	~�e}���gKf��.> >D�t��Wv-;�	�y����B��8����U{#6]����/"}\�f�}��hR��(�̚�w0ye�\�^K�o��-Nk�z�P��F��K'΅��dJ���|@`���V`�&[�
Rw7s��7r��vP��dĺ�Kwa�V��� F:[N���5(��2r��;���fhAa��#�~De�n�?���;
����fU��;@��>I��9�3c"?u��{J�w3rV��+m��)F�i�\�U�@`��MZ�$�l��2X[�-��E�V���⡁/q�ki2 �1�����P_<z\%��<[����
����v��!�h�t�ܐd���S܎`�$Svtkqp�L���e����&�4�1�|ֈ-�v3�db�71;����\ǒHp�zw�3(8�$��Аa���c�B_�w�A�$(���,��׶�hf���})r8�3���f�hu}�~�G7� �7[&^�04�ÆLZP�鄗�[+�Q�G��]?��"�}��u�0L���9�c�{gc�>���3�?�)0�(1u3�� �wsm�7��Z�wb()UA��VNsΈ]��tq�_�g(��j��{x��t�!�WY8�.��G;�����z��|9vo?�p��Fv88ӴFq(��oNNl�*^]��"��޿��nv��"��E��SSm5|"��ĦvT=bv�<���L�i��!1�E����(��]���r�nno�,�Q���g=|�fϧ�؏�U�5�\��0|A׷���YY� ���xVZ�!�@3��;� e�3�ص���Ъc��z�#gi|?O�x��^)�%!6�gO�G�"�n��V�gX��
u�.�v)W�7O�-}�΁ZA?9V����J��rfΩ���B�wqU�?n��F�5jp�it�"y
�fO|�m�R
�Խ�=��������8�Sӕ�0|�er��ዋ��H�u�iJ�X�I���5L-��c�d`�3�2e��^^S�2#�c #n)��"�|�xu��gz{;1�uZ��X��ҭ<_\���)g�D�����@��ո_�)>TA�|��`��L�i+��o�҅����8Xgc�K0��B���컷M�����]��Z��7��Ƙ/�����2$�{B>���ϔ�Бx��/�"���3r��?*�_��Z��e�Eř��� �G����*[�'T������_h�A=�h����������3s
�7�Ӷ�� �\�!4_F��J 	&(6)���K�Ǐ��ْ�Q(F�5᭼�si���g����c����۸�+�'ʗ��^�NpAs�Y�:��Z#E�2m`g3���z��	���P��dMbWCIP�2��Sd�HB���rFnlh�N��]'_��w�טh� ���ݸ�D�B�=�P����\D�E.���`q�2�跴��M�AM�Tp���5�������%�ʪ��C٥#br椊UB� ��a�7/��y9ό�c�zp@Pm�b�/���oT@�ș��55tj[e����%q1V�&�՜���(�����k�rl��}�VٟaAQY>���` �4щʹ��Qr�?���Q\N[¾�(V�� ��,:�o#.�-}bǦ,��,����w-�X��@�t|�E�Y+����]ʬ6�n�w�`={
���R� !��8�'{�����U2\�Bcf��x����������#Q�N �i'�?���ܪT$�	cM��#��h�7f��$8H�B6���\�.������ɒ׽iD���ϯ��Ӊ荃�V��@6d'��v*&��,%��6�9�U%3��*�J5��eȚ�x��[�z�gz;��(��#ܥP�b��C����7��?���q5o(ʹ_����-�V�_X�Q�p�}J������v@�?x����{|���˷wE�S���3S��b�U9�̓Y�P�^Ʀ�&�
�s��n��P�Ow�~1��g2��Z9����,��M�X؞ϚSz�<�Gu%��z��!OMG%r�O*�����;���tߤ����չ���Pu,�����nݡ��r���̈�����2�p(� hP�o��Z�6��r���\bcB���_W�g<��N�3w�ji���{t����Qt��GEv��aVI��1����v�6#�����Y��>�9����ڏP�?��z~{{���������3��������I��@?KL�kǸ3hlrÍe7���ԽM��N��ZY�f��(��l�x�5����.���y%1�G�n�H��J�����
M	��ʛ��&=������
+�+�����.ȓWEjtO��!;jo�i�VO�osC��ʺ�M�\w�?�^6�`Jw�q��J���!z�K>��w6C�XS�HG���ٰ��)�A�XJ�3g�`�������1)w��˒G���ʔ�6��Ė�G�]Q�k"�7,-��o!� p�v��Y�:z�Ae��𩈪��1�/��<��5>Pp�o����!��Υ$A	�L�)j�E[M�1�_\�덌��<�����=eZ�����qB�~^�;O�g���Uwp!J�o��&�k-�#.����r;���ɈtcK��lG�8Xq���5M�YK-���q��̙G�p<A�	��0�{ ��uEZ�/bŗ����*Mͤ22;�w	����k�S K�o�[� M#��� �B�W`f$�z�Q^݅�;95T|��:ŘX��i fZV�n���Ag<���PAiA�]=&��Ɵ�6M�n����Iz��7
RR���O5�ׇ[��$s1����k|����X��_s>FQl�{V9�o$��R�sW#�-Ʋec=��2:�1NT����RD���Ԙ��ٙ\UT1���&P5kX��b+W9��b/�-X9���!}�~}&�
���zMi�8���`����Ф��X\LS��eѸ~���n:�>eT�@� OQZ�
���@0s�?���[�A�괗QS���&~�nD��/��L>[�(��
��1�M|�6FVyA���ݔ��w��X�IO����Ӕ�l�Ϛ}��!����Z	�]�{3,�D �E�c;cn"��&�j���sa���`���?k�q�������@�y�Eg���F����Ќ�Ys��r��efm�h�̭t���<7�6������۔dQ�?:�]VP�W���B�i?������(�>-�p�p=#$�.��ry����j[W�Ī@�C���;>��t��/�(YNz�x���#����Q慄ւ�����\��	�֜��|ǣ�H
B��ɶ���8�O�6b�x�v�f�8���ŧ(3����T�1t��ߠ�fx�Jh�Z���%zc��m6Ӯ�R�C�c�tB��Jz|����������ٝ*7;>��S�īQ^t�Z���oN���,uΗ(ޮ�-�W,��6/<
]����?8��1h�j�L���O׀����,��}@��d�to�5����3=�0���}��i���DUbI�<>b�݇%?��O�"@_����X�;���I/Sݠ�}]y��h�d�x	�ͅ5m;5�����yϱ`�1YV���������|}e�#ۺ��_�D�3�+�mI��zh��˝A�5��Y��o� ��l����7�K�j�������J�.s�5�pQo�DeR��Bc���%����ޟ�����$��U�EM������� w �|'��ʀ�����)Z��N�h�jdi�c��]��χ xZO������:�]��U��J�=5anΐA�ͩ�aB�j���r�s��G)&��D*��2P�C�B��w`�
�Ӯ�2Vk���̆�D}�|��=��Fׯ?��Ա���`8�L���������fs(����33rM2<z)L(S�o���׽���+�w�D�7�<�����CZ�s7Q���)�+%|{��v����mS��,{����O�U��̗���,�z:_H�ꡉty�C��I��OQI)Kh!�:�PU�ʾ hS��֛�n~��%��q���U>D��^����z:�Z ��;}Q�}a1�n��G}튇7D~H�5Xh���x�C�����9��w�v�����.�|�%cr�]�]����>�A>��fD��J�'p�2����O��(�Op���ւ������J-�|SY�zyq��ύ�:�Vx��Y�o����5����6�K����>��{5z'�`p)�L��L����r�u)���R}:��h28��&��'=NJ���ݯ%$��Ba�)�#Ӎ����r!풪%�����K�*������ o+�U�q�0``dw��r�T�lھ�%c��<�]�R9���t��� �G]�R��V�6�+�X�j�nՑ׍����]�њ1�.��͞�p�~oN��y;��>��>�l�GLw�����	'.�ӓF������E|.�kQY�5����d��	�M�ھ�t�c�j��Qi��C�p���J��wO}Ԗ�_j��}��)�_�X͞^MШ����\����./�V�;k{�¾h�g��HDȫ0A��]t��U�2sl"!2䘪�1���
��:N����8|��j.k���'����s�Vw#5?9��u�t|����D'�C�⑺u�h�A(�%�c ;8��1]dTm��hp��e����^���5����9�H�7�wSf�$����@QZZ_���
^v���VO���j�n�7X\r�I�3�݊�sz#���]��P���gc�"���\���n��8�g���?���Eo����J���zv2�:�$��8P�Qyo%������D�Yr��h�-�i�Im�N_��SG��)���'�:���Rhhr�ذ(( �[����	��d��&�7�8���cߩ9�����QH�Q\=��K���d��$pza����s6>����/K���	.���[G �#�c�I�h�%����$��b�3y�+�+�G���Ԃ��$a�r���?^NkeY98ۨ�ŏ�]v�lNLK�d�A��?\�PM�6��ww���Ip'��ݝ�Np����5���K�{���W�Vm�L�>�Ǧ��`�T������(}����b���l�]�N����֜Ϋa&8t�/�I����+ᶾds�����3��[����
��;�;���N���+�̈�R�F��+�jx!�x�o< ĕ�H.Pp� -a��q�>��ۖ`�[�n-ը�,�_�w������;�9sa}�YN���hYٴo�̙9cN����y�/����R 
�ΝT�h����%�m�5T��Ei/��^��<��U�����b������&��~�7�g*X��L�P>��K�I��h��"��z}���_of;<��oC�X�Ar4�9���`jr2�|?��t�P�����|Ůx�mߊhÑ _NF�����\�����z����z'YA2ޥ�u��G1͹�T��R$P���M2u�V��	:}(oc,�R٣�]��a�x�T�B�q�n
9͈@�g�$�ݢu��]��=�����ݚ����T�'WU?���� �ې���.�6���>i�s���4bɚ�z�7��v�U�T" � 3�k(G�Ӿ��&�kn#���Y
��P����h;�w��G�t��� �E�탚)S����?G<���}���e�|�U❗t�	bҎkG�&�U
��<d���`�V<Jb@�%x�k�J�ɼ����A^���;)NH��7ӹl�k��ز.<}
����{� ���Vt�t�ק��󉇟
����_
w7ԾU5ѝvy���H��Ǘ����p腼��N���3� �
�h�X/��tw�4ެڿ��dG4�$k7?��~^t8!�[�L��a�k��"F�����B*0R�,��)Ȑ��Q�u�a��袲PY�R��t�@V 1S��'�(�vZr�L�N��-�o�g�,"�	�e�j��B�ۊ��Sۂ~0@͜�`8�M���>�Ha��E�eTßCg��K�[SA ���'�h�|Z�>8�omwۚL7i&�o��li��mn�z�>L&v(1�ʚ@:�R%�)c����l3��X��rũ���Gk�P���>>�YĦ_��T�@_�F.j9`����^�r@%�Q`��.��ѵ!���+M��\n�c���c&�ˠ^�R�/�$�C�� ��`\�ޣ�{���'��{}�ϐ������\{6�@-���8��|����>�*��������F�5���Ve�h(6ٹ�ĐY�&�@L���8���⨆~�\���.���aC��n�W�B��|26���l�ޞD�����%|>#������ rK�@cGs�x]iN�T6���FA��ɭ��O������E�������dn�ZsjMxV0���]�,Ґ�&����NU_&7a�ݢ��!�&����/�?^.�l�.8}\v���ˠ���ͥ� m��9,�5�Y;�CƦL��|T�#�(�����a��ڈ9<��{�4��eR;�~�);ZT3�ׯb���� �G
�u�3�Ɔ=�u� �r���]�k:�S�y�`�Z2Z�f~�_ێ�h�W���z��,O�Ý��Ew���̳������h�ڿ&�(�eO��gk-*Y!1��ٖ�R*҇F򰴔N
��_'�Y~����K]PR�_�#k�u*K��
yS�?_�f� �2H�x��{9�,"�6��gn����za��Br�)
���M���)�boD�uT�$�T4i�W1DBdt��~if62Ipj�MqB�x	�ټT�\&q�U��4�u�$��..�싮sH���?�AĜ_~I��{�q����V��Y��:r��v3�N�ufÿƒ_?��83Ctns6��=���}��S#�^��,#)fMb6T2��g�euI��Vev1�B�9�Ɵ����%`&ʎ\�Z��-.��,�M�~|���2M%T�1#����3d���g���dc����������Qq�ֹ��pi&!�:�M�r7��1A虌 Ƶ�Ý�����,l�j-���	�P����ǜ��:�Z��͓�<`�"w7�4�_;4n\T��q�yJi�	a(�n�3u�Xn?o��~�M�۝�\!\��jԿWm����}1�Yyk�ܭF�y�E�����Y��r��˟�b�&��(�84�����ZC�ǚ���bӟ�\�`����:���I���M��(_���V/��l2KTT�W�5�@$�(�h�OY���Q�*��J_�C�����MI$`�NDQ�NF�(si�߁Ȱ��,�/�Z���(*2����h��P��°�
��*ۇ�5���C^������@��A����:��q� �!�N��XK�ۅ��	��c�M9 �i!���M=F�mР�a��������Ba�@	��}��p�<��Ŷ���Q
�e�/��� 5ġIa[�cM�\N��
�t �������(?(��Q�/�+��O���0i�'&n�`�bV�]� 6oG�g�oH���l� g���3BE�jq#ږ�����u1�+�1'�p�`���7/��dP:��t�tX?�Qw8�W>�7���K cW���2	�� �Yy�)�q<z�.^�aL�$�G��ԙ�W0R���!@��W�<64���4���(^�Tg�x8�W#���S� d���W"я :M�� �2͹�%��ۄ<tX�x�v�z6�5�� n��$��7�Ǻh57�`h�����v�j�A����q�q3��nY,� ��rc7�jU=A��-:�36y��9�j�Yxy�"q7��0��0��98�����DN���\n�׋��y^T��⁐��)�@�٣�h�����������'�Z�Mqi����P~�N���n��}�9�����@�b�|���rQ��/�fs�qa�ys��L�3F��P�b�[�%{��N�}����z�XY��;��E���{��q���&(��O��MV`FD�޶�{o�2l��xN����x�O�6<�uU��{�����e˟��Ou>'p��}�`9Jiy>=���Z����"!߸����#��D�⿝����m����h1>%�a�ޟ��6�$C;�ھ�� 7P
'8v0m</J�^�W�#'��K�å�X:��o-��Am�5 q1f@�����V���A���Ⅽf� W��'���53V�pX�j[�ǚ�y�H;��(� �!Iwk��4
��ԙ�`bB��}a�����6���]���κ��KM硜�%T��d��u
*k��`ط����Bt�Cy^GlYY�;ᯏ�/oG.O�g�G��N�2��@�'���CG��zn��u͏.ô�]R)�˦�����eca]Q�]�X?��Q��;oJ�.6� Tcr��V�/��t��YU	�Xe��jq��O�ᯞ��yY�0ga����������
�h7QA�Y�-%���!��.7�#�[�\���8�8^P��c۠T�8Ý��d*�T�����ݖ!��\��b�H��}�1^^��U?݆�ubr��`Z_����c��-�m�O�!
�Еￕ*cA�f��QKs'f�[y-�R��> ��Ç	2�U�5�c��~���b��|�)�G�L�����h���-X!�ƒ2n�0{��?$�s���z?'��i�XX]狂��6��e�]�:�.^7�f?lB�p6Z��6(��O�y�)�Ο��f�����p�Ѿ���{��A��Vd�VIvB�%/9i��;鮽t�p�GQ�L���/�)SR5[�������]��Q��S`���S&��뀫����b�5�%�"bMض�Q܁���E���ع��Q���id�!mr�ag}D���X���k��x���?�d�}%�>��"T7�r�A���N���χ�SUG�X~�q�T;�y8xrySD0u��ZG��6}]�=��P�ӳ�+�����;�Dux+	���l_��!
�3������.?W5=+�\�t�6q[��N�9���?�0���v���v?���j��h���j���j�߈�`�W�.stf�/y|�Aq*R�/�'G���9<v��Y��Fi�6�;��&"5;=Н=���_��wژ�	nV�`�'#�O'�VY��߮ZUA�ŌQy|�hu���Z�h�o2����j�N��4�� @��o���&e���'�����}x��b��ꞓ�LPw*^����L�):i���M����;]*�u�$��*3z�7.M�O�ȹS U8Y )2����)O��x�f�E�2+���k��ꔄ^]��ݡE���K�U�&��=� ~J���u���5c���^���ӂJ���6�	����I/<�;+]G�6�Wmq�ko �_s��/��E9���<6NZR'��@ax��ǟEK5Ê�y���dO.������~X�IZď�n��Q����r��;�v�M�{8��͜Ų��1/�K�p����$�痀UY�S��_XL�Ȓ49�zY0����6���F�P$����2��ƛ�QN��Y$/���^l'L�l����^Z�N���	�~
��|#���r!<[ja}|�NV.�ˊ�H��SD���MT�:e�0�O��4&W���]j�^zf>���c�˘������6�( �i�mp#3(��&�O����̈��l)�P����DK�b���
鱃��=��ND�tc>T$��j&{�f4��jB׶�!Kp�����>�Z��v�4sʛ�Zz~ځ:�Y�Q�}��`�|��%�0�9�5���ȷ�d�{Tp�괕j����d�P�.^5]z0#6a�;(xBw�#ͷ&\u"��ڡe�Y��Hg������44�	Z���*I�/�x��%N��傢�w�'����i��	�;�AT^s~�����h�F�Kp��ٸv������GX�%;i�
�ڵ��\ �����]�VP����+��e���l��ͺ�ł�b� �g�
�	m*h����e��sTG&r��-�F�Bĺ%�|5��w��P[�HEJ����ƻzwHU����K�x;�g!�Ì*��ݑ��N���|��h�׬�jB�ྃ���i��3�{q'���o6}��r�,��Q��[jj��*��M�%ԁ�E����� ���C�Ksر5��9Fӻ��He��ޓ��hu�k��bo�͛���|�щ7�.JK�d��N����8����f�H�.�f�B�[/����,Ka(�Bz¯�m5���8ۿY�n�"��&�j]3�k&�b���J�J�W�<Y�%eyI'�3o�$��e�L\�iD1$�}�y����tC>e����k�%:��؇ƴ���_�����ݘ��X>Ƴ��&����r����(��]�^��p����X*�y�.�Ω�q��W�����xE�����W�T"��?��BxT/����d^�x�b�% A	�����`�LA���ب��d��N�DE�\����`��0S�Qf�ƍ�cX��(|���G����U+s��u˾�\F���y7���3WE�]���0�d�gu�M.��J���F�}�J�>��(Y��?=�<��W�����j�ޅ��#�0l~�떜^uPTn��V�
�^��y����]D��o/1���;��Y|���/���I��(q��^��ZGp!/h=��ͬj+�~Z�B�TO�|y�c)Ops��p�%�:�M����%��;��ͫ�L�֔5d�L�������|,|�꩷Fc�!H��/\ډ�7C�̈ǜ��Y���ﱅr��'�ԯ��q�ycl-��?�~2��<���3P��;�whUµYĴ�]E����B�١mM�g+���Wu"�u)l��=Lee�yX9z��##sEY�Lӟ�-���~��54z�c0� z������Ji�����fi������jn��?��$PPz�6t�ĻUO��/����^����׮bMz���ܭ�N���U�fF���i,�.�$�Z��
<�F?�����o��-���}O��퀘嵭�����k�]���6��w��؉��+|^�QCe'M�S�>e2#vі;o��}'c�n�]5�����;1C���^����`�l	T����4mm�؆.mK{
��������I���� �}GHy��r���|9A���N�[
ݳ��8����K��2�e�ڄ�<P�.*�xb�W����Vr���S����]�|k>�r)��Ţ�r�x��.<?̍?��'�x�jƌ��e ����~��I��"�o�H�8.'���۶�����u���c�t�pү�ɐ*��S���;��l�}���lF�+���l�]A��۔�\����۩�_��QVD�������t�Xלs<�/��<�,����Y�~��>xT�����Q��_Oxm/M�����Z����&$����FF�0+�[Nz�7	T�Xv��(X��O�,�3��,=/i����T��xM򺡵XߙTd~-Y~��	��}����uR�
��p�����kl�9�U6�̌x^���-��{>X�Z��Wq4ѸЧ��u�jс���;�E������x��Mh��__
Kz'�,c��wrZ"�`�6�Ƴ7peZ�o�tdeȄ/hkJa�KT~�6�o���7�������ڻ����`�ɿ���J�9������ۅ��۔e1����9-���1���y}�1y-�5����e��e��4���I�C�@��yo�"��G�"��i��O����ҥ\4�ٿָpXN`>�@B/hH3D�.���}r;�5��	��aK��X�Y+ ��*���i1�ݗz�qĮz�8���Tp���n�,��'*�O(T�K\u�
D��%�H4�njuu�֔mU�,r�g۟��Y,��hO�;�B6M_^b�t�g!��;�P��-�z���$�.,>������x*�jzpsD2��T�C���Y:�y��@kUȒ���:��k˹���zd)��ok��t�yW
,.�v���|���ꌐ�����+m[À��*��I����"	�������ލ9�/.;�9R��JӔ�Y㣨�a`+MuyS?|2B�i�9|�K_���XLZe��F����~e�2X)�1mª�b��;����Vg�	]�S8	r�/St��,H��T�e"��-�56W�
��7/��o��[�$�U�(F}\�bL�B���
<B��K!��g���,���-i\� ��!�Jcq�T �w�Ŀ�?�!��\���CCi�Z�,�r�)S�<�����in��P�zw��|�}͈),O6����,�~y0��H������^*���� g
gƑO{2P-����<nЌ�ա������5 Uk���3;GFY$�����7�%!M�h�5�ܗ�5��{LT�*&��Lw�7�&pj�}�ͳ��?�x8�)����-�L����ū���8�j��a�=C�xT+���~� i83J1����)�ҳK� @|��M��I@	�fA��r����S5gHN��z����D��)���0�z
��Q�q*(�D?���~�lV�O��7O�=��K�v[�$����L~�Y�1@D35@}��'��7���? )j����fp��kh��a�Bu��`�<��Iv�����
^>����Kވ򌦗R��1Y�G�T����H�[��Q��~ڵ�d�"�Mh�S�>��cŦ�eE��S7�D��F��+��,�������bie*��?�-�;vw|3�@vO������_�=윲��@��,.=�q�oh���9%I��W�p��w�`�2?��,���^u��.�Bʕ?���n]S�����(�7�G%I��c(�[�Q1�Z��u{{�G�Ν�`[m)(��A̿�&'0��D�����A�+g3O (L����t�V{=����S�d�-,L�h�f���V^�0��V$8�=g�Bt�M�e����?���޳R������>�J�mF����q�Z��n��Q�P6
�<+�{d@ÑF������%�H[�PeW9�'#���]�%�3��c~��&-�S��6�s�A�}9;'�����kr���U����
�0��n71R&��U�TN8����A�ԁ��Y�e<�'��`*�SF��FC.�:e��<��<nd����D����yB��1U�d:�J	�BZ[]>M G��`�z��r�����K�������ҦoW�Ar�m�烱>7p�[��X}����R1��0D~kU
c�C��Y+�����l_M$�Yw4:֙�5��)�Z���A��21c(�`�V�I�5�K^�%�6|��P(S�q�}�-�h6UУ%/G��b6�o���B�z�WA�����&����x�|]�\:��C��Y���ڣ�v�R�B�}k �����:B9Q�C#�v�LnP97K
���ڐ'���	��H� �XL�i�ao��!��}z�,�GK�=��:��3�� �['T��I��
����i�ې���1���PDq'w�@t��1���	����O����Q_�
��%<8��1q͌a�g[�#ƀ�X��ԧ����tE.XCW2��/w2���d_�"E���|�EeNg� �D�ŽD\���]t�!�������]J��Э�j9��u�CK�]��|����
6J��}�m�$-��m�yM%uBT(��6Mtn{܃�XZw�7?���i��)�֎/wBx�p޺�0H-4I��b2�kOI��/�N*\��?���Ew�NB $�`�-Q-�����f��c'j��O�r�+�U�3sj��zT#�5٪�P��Ũ�Å��S��v���*_܎����AN�P3�����l�%ku�]=_;��$�
���z �A�Cn45�� �ǃ�|#*�����J@Ir�O�"��Z�Ѳ���dKC�I某�%�p/|�žJc�L|?u!�� 7�j�	B{Wx>S&g�ɟ��1��#{w�2�c2�-���(�Yy�_X��s����t�jL����0$(�0���5?^4x�M��J��j�})}=cH���kCdK$�-w"�	r�ñv�]j[Bb/�z��Vg̲���8�L�ispk�¦n�L�8)�����h���J ʅ�4��")H�eHX��l��m����L�e������Ӻ�s0��������7�\�B7��
F�C*hރ�����PCg�����]3(����ǉ��8��r2�ڕ�B��bV���6DT�/�=�+�V&NV��@���w��.� �C�Nn��Pִ�b���=L�sZv&����@����C���݉E��d�g?*����"z�K��xg�Î�%��T݅��Ϣ�~ ܎1�/��s�4��ٺ#n��\�G��W.���߱�"��e&'@�Y�Gf'F+�����0������(�gr9�T�Gm�;�{�fG.c�\�N�"j�nn�%!f�������2T3�!0�8��=���Ϛ#tbq58О9c,"5QqbA�S_4'D�M�{!���>�#�8Z�rWn6�<3�]��{��Gf�;|�b���'Fڷ��CB�%���Ɇ�5ﵵ�y��υ�De!n�J#�~��%P�D5��o�� ����g�,f��Qq�Z�t�_��d*���EX8��KhN���K=
\Ծ/s#��#ip^?�������B�G ��(���:xܕ`�:`:v�.��A.��_+S\�a)<�Q��Ԅ��\CG/�}�ق��9�Wf�)"L��� ܲ�X��/��*%TޝZq�߱
@�dq�?ŗm���#��@<�Z��k�kw�g�I(��4>[mݱ����%anY�r}V�V٧���K��@���U�����C��]
D3E��7��T���V���2GBԎ��[86�A�V���..�n�������x�S {-�DG,2��VM�| Mu&����*ȑ��H}�u�n���=&ꐂD�@��ba�K�M"�?a�S���P����0�v�)�w�l)	��a��)�0���u�����K����9�ޮ?|:��U}�x8��}N)���_����D��$��c�|�vzp/��j>��o�[*7R�*�5rT0ᴝ�.�?믔���3V�*����%8VUJ����f���9"�oz�s3m�j���� �{�����������	nI,G���98��fG ,��;�AgMP�=��U��<R'���!�Aȫ�SZv̩�ԔI���1`�l�~h-@s|��R�N�j �C
S�tW ��h�oD��D�=�m�����xz�gơF�"}�G�z��A�|6���R��ۺ�O �wEۘ��_�����i�n PL�&���R�^�=��?�*j~@"	0�UV�WB�6ħ}+����)�b_8�6�� \r���>��v����,y��%'n�W��z(kh@(��ť]�{�'��g��I��j<A		}����`�u�S��Mn3����s��&�E05MӰS#�F#�YLxdi�i�s�#�w�|z�0�&7�NPA�5Žߤ�����qy��k��}������2UtV�J���֣V�d�U6������˔������.���2�Ƕ#7�c��EO!ӛnlkty��k@`]�q�d2fF��(}����ʡWxu��O���EjyӃ�|
���R�P�%o'�Eܝ���}��{v��1a���}��P���(�W�Կ�۪�Ѝ�ܖsmM�q����$��V}�Z����c���Ыv��P���\(q�L�W��U;/Kq}�����vb��#���3ި�Y$A����+�U�򜣆�����P��7j+���Z`*?G]�;�V�!%�{p�ޭc�]AA1*�ڍ�op�՛��+����!7xD�<�w1޵�p��K��z�����.0
=�7&{H��n��IS��s���=/g۽r��8���������.vC�и#�	���+[�=��jqC��(�#3:�aB�B�����Vj&����6��^&QM�T�ϥ"b����Yg1T5T�Ŕ8XO�EP��m��b��r�)O	6��X!����A\Y�6�f�(��k�Y�a�oY��"�M�X~�Z!���}�w�	n�V'��� �r\��Z7����vzƴ)!��6��aN�L�N��zI~�����z��ٯ�ub���fDaBX��;C�@���-�f�^sbw�ۇS[,�ޚ!-%��5O$����,j�y��#Pn����#��0�K�$�Go]n�]gi�}o �*4�ܟ�I���S���c�88�]�4���L��	��?�|)B�q��*5Ǝ���b �JUR`���]]�7��[_Β��!�)��4��������w�s���*8���m�b9����������K��W��kl�ڞ��=�ia�X����tfkjB������u�����y2L��cߣ�uZ��'i�e҃�r���f�~K��a}��5(��H�����w�3���!�H#2?L�&T��rw�p�Q��LBB8PKݤ�L#��
�Bf}�Y���˷��A|1�4�mw��w�:ѷD�g��͑�.7�������Kn/Ab���a��)5J\P%8e��c�d닯@�.�2 �]���8g4n=N(J��\�]s$\|I�<��B����\J���"G0�ln։v18���s&�^��������ڄ� Ot9w"9n��苽���c�Oޚ���Cu� c�v�B8&B�0!ב9��~��^��_�q�Z9�ü�6HY�2Z�Z8��:,'м�q4�d������)z�"���W^��C��(������o_[��E3�uiב�k���A>B���v�R����i��Җ�װ}�6~���u�����:�OG8cwtQ��\�T={ʬ���>���D?����3Ӳ�:A/+�q���֭j�\���a�t�n�z
�L��Fi��O����kԃ����������AL�E������nO�ܑ=��ҕ���u݆`����,��yǝh�G���:P$H�T�,��hr	��>P1�j���тe(���F�x)��x-�N�{��~R� @K$�sR0�MJ�8�ǆ�@7e��c�"��LØ� �.�k����@��Y9�&%@����w����:��S������]Xkt�Xl��:"�<�<�z���}�vdd:��nl�Om��2�v�E����<����eGh�u)Ռ�����n����R�w-�w�%��RJ�䲥\�|���x�W_u���o�;W�4��� ˃� (���	��ghG��@�]P�����z�2�8=��xyW�?�R<95�[�+ڋ����_��s���q�}z4q� X	��5TP���������	�q���F��1����K�+	A�q������͛�0S��1C@���5^9�T#��ۇ$���!���3���s���8tn:�v�k����˴r"��ͧ���ϊy%;��,���ozB��D1n:K�L���N����b�q����-Y�EP�#��1w�=O��Of�u+)���n����ǎ8�=����_S��r����,�Ӳ.��:Oڝ�m���F�I,c�@�|�$4%I�����`U1���׻t��|�ھ+�̥=�@&<2��v�/:���| ����^�3����; ]ͪ��<�b����3���^�����xL�`d�r��c:�9Wg9ƥ��FQ��M�	NB��~+�����ig�;�-Sj&��^�x�}n2(���=;�(�v�%^o��X�$����S��=��7��@.ݜ��RL���m�jG+z ��i�Х�$\�B7����s�@���5�׌��|3��G����,���>R�^����ł�A�*gh;�S�iP>�KCy\3��q�Y �2��T�@��}�a_�!ۛ�t/��<�ܝ�:滄s
iLn5��-5��FP�v#�HN�I� �����Vxw��i�`��²<�'�+��m�EÚB�<9b�ऑ�c����`yW��"/���$�β�Z<v��.�mVX��A%!REk�n@2�Ab"A�#�<��2^�^[��d ���O������ڸQĶ�UΛ��	���p�ݼv��������0����B+���F9Ll�8L�6����#32��oU_A�
�w�1�m�04$��;�篞v�GP �'V|3rp�����^�*��16�_�!����5�%�t���+~",���pQ�g3�ytE�E�"'�\�Ѹ#�A��qю6dJ��K؜Y�-LTgꧣ��)j�Q�/㱣f��}�
�_�o�z��ۘG
�u�dĹ�β���bێ��wo�Ce+�O#�������>�͍�Y+Z@�nB��$yL�-�FM��|��D>@�F�O���bW�ڔ�g��)�.[�ZF�.��7nù
��|%�p��9�vz�>���V7ӵ$��t�������ɀ���ψ���2y7MY�!�((����'�曅 �����t�����y���eE� 9����*>�R�M.�-�B#Kа��i��d�y*�Đj�b$���
���|3aF��G�l8��@�{j��z&X*� ��[9��P��
��~/�/��<�� HL���W�9X����<P�P�������.q��G@�I�jr\���|���n��j��?��1�V'}�C
�C@�1=��06��
����W�v*e�;҂з��-pr�i�;�o5��ey}���-�>@T�k�p����
����V?�ّ����124A��ڣ7y�ە	��c` T	3&��!��G�#��p<���P�������M}Iq $���f�*�6C$-����O��`�OܜI�vyk��tc��+��ܸ�X�v�����+�ҒR}A���1,�8'����T��?(�~Z_K�j�����X	p;
k �>�ǕږlL��0�j;���Q[8����G�2������ S��NAVR�<�����
����y�7n�5c��+W4<��b�ٌ�=mK� ��0�ҴЂ��BR���_�T��>б�a�X��Qg�괔���Db�K�@<3l���6T����YQ�2	��g��ĥ��K
���v:�g:~����j�l5�>C5�ﳬ�����oij��Rl�l�i�p�y��L����^���}�L���d�Ӏ<7~��b�<Y���t�xT
��uC-�Y:y�QT�<�X�`��7/�L��d�?�GXL�|f	p���P��m���z�7�VfҸ�b�=���c���`_��xr��H�po�+l���i���ޚ���XH=�C�_t��D�cP����.�BMM�J�����aO���,3�+
��7YW�F0L4gn��;��
c
n-0*��xTC3	f���I�x �=m��\�|�� l&J���/v������֗������>�a��/���2��A���jВ��
~ �F�8��h~�C>8mu�a���t�Y~Q�q8nPq��A���	�G���A�hŊ91��;�����~(���:F[���^ۯ�A(*~��CЁ`3��3-����u�Et��kA���I:�C�wE@��m�vaiv��:gv<	�vFu���8k;�ݹF�u��c���GV�iJ��v��a�e��?��aM���0��ޛ���iV����
�zh�U���SUQ�5���b8�P���Ga�l��@菕��=�a�T]=��r���3awww��f�g���;�Ƣ����:������b�>3����g,n�hʆ<nԇ;ԉ�;����q���/	2�̰P9^���5�Y��A<� ���wA�,���6����/�74>O39�5��0$^|ߨ�y)>o���E���f�'��ۨ�bZ�h��C���{r��P�� ���b�yl��{�^�� >��7�ׅ�����f��qes�G%p��mGp �6v�TYY��M�������dw��|J�!')��|�zP[�����d��/)y�诣���DE�_F��R6~:����`���CU�m�Ŀx��.O�'��B���>J�]�]<�ĖO��J�	��f�kJ�E;�i�� 	�W��B/��D_�x�.Z�km7��۵��rVI���\U`�(�O���|�[��/6EV=�+��v��%���ܢ8`L�+�#BR�1zZ �"T�I~q��8!�5V��pi��38q��T�Z��Dr)���Q���s���܃�+m^\yt-×�lT�ч�3�|ot8ZR5�bn	2�%`��04�d�aB^4��{���U�T�Y�,�E�S�P?�/G�&��iq���j��	C$H�!*��s?P2Wr2vr�n3��C��SX���A�ik��F0�R�� ���)����G�Oh͑b�&��k��ς��E���Hg��H8
O��Y��a@��� ��j���C` �B��TJ�%��I���$�q�Oh�K
���?!��Nh�?�B�����{��܅d��Z��-
+#q �y�s�Phm���a)�`?��y�?��OB�lSޏ���s�&*}�5t�w��"��?�AS$�!���|�i������[D�jw����?6���UW�̟���k�L�`�����CR�[42h�h���Cⶅ?�R��2�5$��!3����ꚊH��G��(&�&��j�'f�)#K�-�&!���B��p�8P�~l�����~� u�"r��\�ȝ���z�B��7��JU	���5'�v�[ag��ߠ����
Q� �A�4�R�!'i�Qg�p�� Ɏԇz�N`i��Y�d�Kի�Iq'�P���M��Wq5�EC�P ����H�
�C/Ifx9�ǒ,V?@���=�?J-�\�>ް"�b�'� ���5�(���c=)zڪߢs�A�̜t�(XQ�4H�Ұ�����2��-� �=DtRf60K������#�}H
�M]i�/��|���߫�������n]iW�}�	_��t���,l��b�= c�+/L��0�!,K�� �� �H*��hPj����J_���s����M:�&ް�[0��A�x ů��6V�ǩ�7���Ö;�o/ w��/2��#�#��)����%W:��$5I1��(j�!���Q�@��$�u=��?���j����u����\l �o���l�+�
������T1�� ���ΰ���Z��[���_]�v���o�3��z���(*�@�L]%a7vR��*�;���7K;��}�ӹ��~)�R�c��[�W�WB�4[f�'��*QE�q�[�(wȮ���#�ז=�������v�7��TV�����:@�����(df��ޔ��Y{���๸~��p�z�y��+�avG�4�U���!��-����j�]��dg�>�B�Sbu�=>ڠ�>\��j1PY}���2u��;#u�쑞��<�:�x���q�:���l�Wj%R�{x[�^�ȃ�A�n�Dl�|��<��%O��\��u���6I���8$!��L�J�щ����u�_����o�}#<}}& )G�òT�H�q����ڞ��|2R�]�3�!��|����g����(Dc���!�	��q�ߗ�h���N�t�/�'�����EB�� �I�����&�T�5�(f���P��"�B4Ht��P�:25��ȅj�#�M�~�^��ܱ(��NC*��N-S5�&����;�m�������f��[w.�~~p�(�����ŏ�����3��A�;l�x�{Ux�zg�\ʱ�%�g ���}�O6��B���M_�?Q�������[t0
����PT4a�hڔ���������oF�2rrv�ԛ�㯅^�q���Ǔ�����j��ڼ	��t�HE�ނҫ�J��(@jD�H(]@�H��.U�-�*z��]��7�f��53��䞳���쳟��uW��E<��J%�И����rC%6dA��{�f��1�E�5m���_ד��Y�7�����)��B]g�O�b/��)���yy�&�4bƋ~U�Hs��uE��inl(���L�jt��`��N��ht��n�P����W���a�雥w�~�JV:���m;%�mB"���R ��{=߾�,���r����7����c�V�,kC�rw(*�e���#���v�F֜�
���^	��g�?:bu��;&Ism�U�f�Tf�fZ|�]ay X�3����>���޹���Ns<�H�d�@�m�s��Ϻ>���|�~���i�5%�s�hc�k?T�v���eH�N\�0ְ�[�im������6L�!�$,Z��ɋ�f�V06}��S	��3�,�q',���:��jģ��#���J��?j>3��_B��t��*�h1{�yI	���T�ߏ��2�kJ�"�\O������_�81r�k>=X}�C�)��>J\g�	H-2L��#�`�V�IǟCIqd����!��6����x�X1�8�*���1�dE� ���^���X�J�"��p-�N^��*��%l�_��ʇeo�^�to2<�����uRVs����\�[qO���m�̗��>>2ҿ���P�g>�&�(�_���d�/�Y��0ik	g���)�
<<c���A᎟-��L�����_{��tv�����;�/R%{��^��ף>�U��W�,���"�3d�{�²�?,9�5�Ɏ��
�O��̴�&j�[/�J~���ݏd�-2"�ʌL��#���X\��~�M�W�-r�#࣏Qq���VT"զ���d���h�R9@R���ё��ExDu�u�?�ѠN��9f-''��>�6��Bt z��ӫ�(�
��틮Y�AKE���.���鞲֡��@k�U?V�Zd1�2�$wW�-d�@&�A�\���A���hSI'T��C�x����&�NN������IE4V��J��JD�Pxj�7�8�^[�t���%:��!Q;NO����;��@��X�FQ {�-�w]p8ִ"�f��[mS�jW�l��Y��#��4O�����j��
��g^T�s�Ʋr�u0��7�\�Օs?|��u��������f5�Qt�E���OP^O+TY�k{~4�|
�#㝬��M����p~��HT�e�_��V4����'��g\N���J�|��do���*pNnnL'038GR㆖�s��o������������+/(Rh��z��Z67_21���6��5X�̙�݁�#�y�@D���P1���@���� ���%��a�D	Gwd�EX�)�1�/SMw;�>��Ԋ���=LS��[��P+ d�95� ����Ŭ��z�k�U9'�0KY�hW �Z).Z_��?�h-�D
�BRr��L���q���n:G˦*"���
XSu���%�����nB����o������_�#Da>�A����(h��e��J\,��E��"�ח�>0+��o �#�[�q��B9�Z������ 0䥮W�*�!����;Z��@�:�O�@P�m��y�0� l�#�/�0U�DH�Y�E�_t.#?T{Z�V�L֗��9�1*��;i�0�m�����'�̽�<v�T�ޢ���/4Є�Z���J��Vkf9����FI�T�ԙ]Q�0B��N���{!�6q�vƻ�
��O��C�R8�����Z�	�Hۗ�u|����"BZ頚r��i�v����ɩ�&���`��:c���mK�0 �},��ϖ�8m�|����a�ʳ�'q��$�W�RG2��&���;�|}��� ����r6��J �X�2$�����R<���!V�a��PI���{M�Fu�٫�04��+�\��7� �_Ri����*u����'�Y�,���"�Yp��p~��6vvvi))���S6�2>Lm�w�2���)����2�2R����<S'H�T�d�
lsC5�4��?<�6���`?+�4�(X_�[�l�k�iZq�Jz�V;!z&�+�����m-�2Rl=a����𺵦'S��9R��btuQ�t��9�/u|"lgR'�Z���_�±�+V�8�D�h%\W��乚&�7�mJ$���;#y��O�z^x_ 8��y{���ADa������.��x=���D_��*+T���07�5e:��>N��(�][�˾8��ୗ;D��0�����Y�8����[�˞9�����q��G���b�ǡ��2t6�<т��`����x���v�>R)�k����'���/����#d={��m�Y	~�b#t�h,��.NK�V�+y�YC��.w�NYT�kI��>��E�)�-�gJ�.Q��B:BHG7��n�s�����/^�s�].��;�@�Ҳ��g����Lwr�H}	�1�� 9fC
}@5�}��i^C�^�V���q�#�9�U��a��~�O?�
jw���\��&%��z�	�`�$' u��:�k.^�׹��{��>�_wڦ#*���_��g-Q~Q�2��E������z�m������"�$�S�|�E?�h\���1�z*���.�c]?\]s:k�J�/,P���S3�_�����_�ƪrEB��K��}&sR� )i�Fx-q��N=D����!AEت�il5�Fh�=�[͜/`�k®�xX
���7�0c>-�{��L���[��m;s�S���RHŠYg{�۷��0�������t?�6�n ���X5U����&���n<��u�r�JH3ou�˭wM��r��%<=+7�C�ۮ�Q����rj��T�|��Y)�N���*z���Wz��Ol�}�~6��W�L�2�{����j���(�d�HY0N� ����C�ng"�Ķ��iХ����j*��ZFfl�	�C_��n��A�6�"$5��!�K�1�z��)�;z%�^qj����b�w=��d�W9]��<N��.�,Y�?N�n.������O�"��3�fl�B����.�2*$���T�g̕/�v_J��?�jI,[e��{w-kǿ�p`���t��H�ÖN�p�m�g9܂-F��2��8�b�M��� �ꛗb���չW�'5ԛ�NW�P�̖y��&j����p�7��p85���[r��$8�֔~0NC���H��k쫇a|�yee�1����'F�]+"�x#��zJir��b�u�CS@06��4u�*Y+�	.��'��ƦE�VO����^]�*C�{2#cS<X�Ɔ�j����w&s���Vz��eE�R6X��F5�g�BU�t)۔}��0{�)�&p�,WEP�tɧ���MV$�΍�2u�8�������\��;�1��𫡌f�J� =�ɒ��w3���W;�M�b�*)��H��W~�V�I�5�O�{���;qx��o��P��锃"����	�A���Ch��*�w�Zݭ�^�O\��dx�i5�;ٛo�ہ�q_����Ę�N{�;���h�W.V0�x��"�v*��ʹO�5n�������Y��	/Y,��7���ke��A��ƎW�]�7��/��)f�Z�X	��ɭ��5�"�j����Ki��fY2D5�ۯTm<v��&=ӝA�m����cU���y#�c��8�O{�^w $��l{�@Hh��0�o�k>و~����2gH+[YY=m!��}n��m�7��F[6�D
�Gp�k�/�Z����ܳ��YJr���8U����rwj�b=cyw�i�����qc�˾��?Dpu2��JC��M.��ޭcA惱�ic0_����+�_���b\g6��:_SC.�,���!Q�]''��i�#��n����>i%���L�%-A4�����V^'L��<"\��saw탹��_��>/,^Y`�:��069���Zu�5;[AA��<X�#:��<s�������#c�����W^R���~uV%�O!
�j��K]$�>i�d�U?z^�����Y=�[N�RP�?ٞ���޾�>:�w�Jq�i��	�\b�����������[bbLKU`1`�v��[��z�ּ��\���N3�f�������sۛ����k��V�_(���N�a/i�~mZ��^h�x ���;�7�[��(�4���s�����M�;�g>n���舎�6��(�0���Q,>�/l�HP��!��3ȁ��� 1��}�Oӕ������L�Sp�w��چΩ��HK��r~�_��{tyZ�`�5f���Kw,�(��<C-�ߺ��.:�Ye̲C����D��$Q]^Y1��(�r���Jng��m�"�5�������ۘ�W0�Ǆ��{���_cA��G��xm��g��M{�n��o�6m��ķǊ�o�$�:e~�.6m�k�8f��g�����T��"�U�&�I7,��t��M�n��C�񍤢߷��'���ȘE(���}���jK3L�rk���A��D@���ag�<eD::J�9.]z���%W�֒�O�H�̘�1餛a;�^����5*�W�I'����JR#9�@W86��tz1�B��!��H�9:.�R�`�+���n���L��r8>"G�!��Ǐ2����F�`]�]gQ�4����ɻk�$��o۟X����{�L���./��~���ߙl
�%�������?8`D
l�I։���Yg�8�����RF��U�8�ň���{M�z�6y�vZ��b�X��;e:)I���?=��o���eⳁ��3(�Ţ�$��{��K,W��fw�d���v��@���g�B�s�㙂�tl<QT@;�~7gw�������V����;�� ���lHK���,�TΘ��f, m������,�=f��y����	�I�m����ӂ��Cb��	\?��E����_��ֿ��.{��������Pq/5.�����Z-G?EQ�	1�%�@ �0�):~�w��d�h��#f��Y��4���<fox�D������b�V�"E������&o�E���jT�b\Z������r�]32���E��-�BCp�������&�E<Id}���"Ƴ���6lT��K�z�ļ���;�4�7n\|��[�J�lp���!�AD�x��0Τ/K��歭�­:�8�+]���ɼ���J�Q 2��]��~��
�)���x�`��D�00��8���/p��^��q�ڲNu��[��{-�2��E�j��y��U�J$<+ #�VW=�q�&�Z��Y �6[�{U.Hd����%kve1���.�,z^������%�'���O��7c���H�+��·}��㶞
��ށ˖hj�ӄ#��.o֯tZR|�k�/��)#y�f��'�H@fXs��n�Ш"V��m��*�U�ٌ�~�p',����~:�\?��P���������\+p�gkP���
@�Z	��;��Ջ���@(����d::���)�R/�v��F�6m'\ھGt�q\���3�;��~�0�Dt�ot��t�ԁ���ͯ��q�r�p�M�H�g��d�~���Jf�/#/���a��ebhg;.�N��r��͠���p��޻�$.ζ��NR0\;�hbi�>��T['B���Є"�6!M�SS`��~�(����z(̋�)�Q����D,7G����`���o��JUN�GƦ��`;S�/XOqY|=gr-ѻ�N��!!*qz5�^k��9ĩ[#3(Ʉ[�8�����?b��K�<Q�$Ԟ:B�n��2�Mv�y����c%R�nL�y
�5Z��w�/菑��!/�7*y0���*�:�]������rtŚh$��ܸ�I`N
�K�n֍�t{ᒧ�e2�����K6NrzM;@�-*��ǭb`y�^�G_��[�_�7jj��1B��c���N0�V	���b/A%^9���y	�r�}`�t�w!�C&�|L�y����ߕ*Я:j�O�@0rF������(��R$�dg���x��S�A>���ڄ��y��������:Ij�ih���c���:hJ��Dm��G\���3�=�F��?b�����������Q��d7:XxCj���9N������(�H�-�%���?x�S��^���< eK��q3�%�e�(+��P>=zs�E�7Y������,�P��P�Y�*��2J�~��DaT�=Yb�m�ű��������� �(6Q«�י?�싴yް�[�˒Q��<ojoh���P���o,����!x��E��k�o1s�n���m�&ry��;s�KZ��"P׶���2UK�7,��.�~�&˫�I qs�QOV�����)�F������;���51���[�G�������6��Џ?��i�W�~/��%������~�,�6pus���fY�	:"�jl�7���7ǈͻ��G�������.���ً���<����`ff@�����!�G[!��� �t�lοi�إ��C�8e�6��g+G "�� N��W��d ��i 0 `M���i�E����n�mԄ .g���w�e�� � ��u����3 �\�Nˑ!�/{ĭ3S@3/�T�T�~������`�E0fi�ׁ�~�гF�6ZV ����|h��xuۙ��; x?S�n�O+d�%hX(�U �
=��]�A���b�
���W���+��
`y��%7�؉������"H��\���V_pOCf���JNoK�!��ED�Q��2�j��z��w�h�|��O�ue�և·�=?[�UC�R�r�=�a��+�.'

�Oߧ�A�>�������+&�����D�C�+1�\֩%�������ww�G���G>���_og���������;��D�큸����������޳����U�n?�/PK   T��Z�'k�  �  /   images/94f8244f-e118-4f93-ab30-835e0ca4f6e9.png��PNG

   IHDR   d   &   2r>3   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��[	�U��j{���zI��t0i�D���H$��3g<zt	G��AFe���(*3"�":.�
!,*[�$d![�ٺ�I��o����ߪ��@:�%��Mn���������zo��{r:�P$�����Jv�W��!�6Uuį��뚃�I�Op~�/���$�v�a�Pw��6�>j/��n���G�6�Tt��}l�St��~�S�J8���'����ċcÊ��h:��<���c�$�	�4@��}WM-M;0��Ј(��n�D�:��朵$��x���D����!G��t?���k�~�����]r��4�4��5��&E�NxO��i��}��\<�a&�9B�o�؈Ӹ�>�3+��ry�]T���C�ُ�ˏ@J�ìkA�e��(�϶��Έhϵ��3!��ܹ�!U�Ba�]�p!M�͜�'�Po!�8�I��sm���}瘊K��de��`?Sk�����^����i��P�"���b���LD�	��0/��ٔ��LB��:~b��*4��t����9�ae��"�K)Lȸ��t�y�GE[�e�I�Nc�W~d�⿎L}�B䉯���\a�d��V���5lL��1P]8
&]h$~�]�,��D���Wqd���t�p����1��jS�_[!b�tϣ X��B���cR�Z`�<X����2Ix��<ԧ,B�$1g�x��qV�.^��H������'N��B>�X�Dm}Y�ܰ�w�G�'f�y��h�2�r9H�	��gM��[�K_�aȧ��R�	է�fT(H��4 �^�&��P�j(Z
REx6TG�9LL1�z�RqZz4��A��"���jנ�	�W��U.P��m�ϩ��% W���ʑC�,&�� ��n#�D�j�Y��r�n����{�}�,`�@�f��I�|#̴i-T3n\>��щ�΀E�i�w$��� fϞ�k�����'.f���2A��A���~F0�'oCJ���(�Ť����j�Ѯ���h�v2�A�tt7��ۢ5I�+��>���� l^�;mC���v
%Ocڇ�N�!=z%�1���DL�����S�v���(�l�EA*�&��{;��ͨ8�MN:1t��P
�;��D� �?C�Waeft�Ǖ4�E��cČx@#f88�ȣ�&���iHU�h?�O?�$�.\H�I��4�2\��p` �H9�~�s;��/����a����0SK�*�a}V�g�F��b����&b�Al���j���A���o���	�]���VPtG�_~Ӆ�k�m���Q��`�ԃ�R��k����ކl�h���|F�5�����=�8O7����G�M����.�@�������G��Ryt&Iw؄h$	��":�%�>�Ïko��h�Q�1��H]y;ꪪn���K�޽�q0��Uo�`�RF����V�H�J�O�IT���Q�OP���$��"�
�L�k)/۵�8��6�I`ŭ�G����q8w��;y�y�������0=��D^��C��/K.,��E���4�T	�����]�<u�.���!��XJ��������7L̲ϙ�2����/���3���Y���1�"�L���%?_؞S&`�'��z�ʛl����9q,�"�d|�T	ӟ��4>��@���z�ۻ�%��!�m�w�Hr��A���+��@:�����A|���&�g����_��IÞ���u�1�y]���e�#PN"!�Q=�?��*b��;���j��i��Sf�R���F���,�aS0l��q��ڎ")(ɒ).��֧���p�Dmď�����t�CUdl>�Ep����i��5k��U��/�sd0��cv}�����m��xlk~E�wT��!̌A;�����R�o�pѠ�|-�WJ�xӨƄ�$:���H��X ym�E�R@��"����k$�:s y����1��fƺ]�8�>&^k�ϒ�G�X+�j���}�\��1�9g�^�eTo�z�`��}fnH������[qo�u���7&p��,_�4!E!�@���-˂��0MS<�w��4���4#&�>g�ْL1��]d35W"G��5̫���v�k*���֭_�K�/G�$���(b�`��T^����ά��C�;C�R�׆��Л"�9�Ag&���B��d�������4MS!Z]�444�
݋��ATWWc�̙hmmEKK��$:::��da|r��Wa�Q(`�h��Z��[�$DolCb������"�Yd�.��PY7�v*++a��0�����Khj�~�k�-|{;��e1C2��!L�

�V�x�Ј#VD0��e�SIn���V���)��kjj�`��Fz��؈T*�={���`�����*��ӧOǆ#q����c�k����y�SEL�H]&�%�m�=C͋������'��ޡ!��ރ��[a�*q�3����%��U����i��r</���l�\�.�ڱ
�)*&�E�ߧɱ:b5��:�Ţ`��g���+W
	:t������/b���طo���3Y\gFB-Y��&���M�@��*�dڞ>pS8�HӸ��B���a�����+?F�#�@	�g��N? 
&���h�˒</�k�M�;�I�ò��Ff!6Oɴ�
�^�7n��ȑ#BE]v�eصkv�܉ٳgU�u�Vq��ö�L[&~%<�� �-%�7�I"��Y��
I��
RY��W![�`���~�0�n���/aْ%�����˪��W���"����'�"�����F����Q�|j���N��Z�C���ǠdNڊ0CX-����Lٿ��f�Ē��mmm�%����=y�5Va����TY *Ո�
�j?yTgTI9�.�>2��:��[!�Ůh9��9�%��S�e-�z3�;<�� ���ݨ�6�*�Y �J���͛�x<���.tww�w�Vx��ѯ������8�3|4�O`*���0� �xW'�ɡfV�D�qp ���]��KR���6m:ló��a��������J�A��]/���"�ߎm c6��1���3��[UU%ο��jkk�!����bH$B���L{Y\�Btb�b�؅̈����	l��p2��$��E��� ��]���[��d%2��E���Q[Uq�/�o.�UV��@-_0����w�<<Sh&�0���l?]ac�c�aJd�ذ�
c;�##W�=X���0q�3���H�H*~��p�]����ds"�ۆV��ae�b [Q:k!�W}�?܃�tF��H_rl9���L���{�xte݄w�F�xU'��J�H�H8n�$�P��]��e�a/�$�y��R�2
KP]��Ϲ��zT$��y����Z�.���B!�-"g��/=$vk������G���éK9!�(/�=OpM�-��:VaO���,I�>	/�\Ċ��w�Q�Q��R��Ҕt���έ�A.o_�("���_{����}��f�~UxY%o?Čס>�?�{�~Z/���q��[��!��ea�Y�k��7L�QJd[.ֻpsh7μy����E��f(}�1¦,$r%�0�"�sk�¸�����J�w���.���_}��H]/k��4��T׌�6��؏.+�K��g����'��#��c���y�`{ ?�R�_T��X$5ў�(�.��l�Ķ�j�^�C[_��T=�����5/\��������tF}Rz��^� ������G���<E���L6V�L�퓧������;}-^'f�j�Ϛ �����EBIlPu�d�He�����8�)�𲊤�T�!�����?q�w ���#b�4�}b?$������p�|Z�P����8ht������K�N�ca���$�r�֏���<�t��,bjysJ<#��k8r�LT�,�h���y�}���Q,oCJ�_>4a{G�n [Qj�;�V�A�{�&�
U#���Zɡ\�����ק�e��gޫ�]C#�a�E���ӝi䟸��xj��` U<=b�;��7��[����f��:-���D�������8���i�i������.���7�v�rkx'��y�	xp�e=7	/��H}��I�v#u���҈؆��_T�lV�8���b/�S��i�dJ�ѕB`�;E|���t�b�e�q|Au�b�w0��f�3T��e$��׬���c΋#�s�nO������%�І^����\�d{!��Mqa�_h��u����"�4U�9�B)ً��F\r�%�'��
��kXa�&0�OQ]Hu�H.�=�c�əʹ�*���O���"����u����1(�%�"ͺ�3!�&�� ��V�~�Ex]i[��i.�[_���ދ�+V`��,�C��s0w��7�r�8O.2QC�	��/k��/�,sl���-�.X��Mq3�
�K�HNID�?�^>8(��_U����3�\9H�D��k��{�݇������-!�`(�_�����.��D�����J*k�)TV�038U���������,�����Nz۽�%�G���f�7�D��؉eq"��� ��N�6g{�,�Y#�!�Oo�}�ń�Kj��a��hy��]E#��}�uw�c�j[���_ �ę�4T�\�=uB�M8>l(5��%�&v�!�:�?�;�fy[Z�3�%�ENw�?�ݬ.80s�|���{~/G�!�a�����
Q��;q����#��A2�<�1Ln��a����,�8�p�p`J&���?��B�``�t]߲C'��v�Z�>D����ؒv�~X/ݏ�?܁���U������xO.�b��)J5ᛄ�§6>(����	o�q|�y�J��~��(8VKK���و�l,F3��S���.��	}��, ,i|�y��y��!�N�sv�z�"�N��&��k���l���a���z��#gaQ�ii� ���K�����6ࠀ�IZ!�#�l?����1��L�$�RQ��qR>>�ʛ#g�X���:1�[��&>�j��Hö�h~
2�e%&�e����P)��u�Øla���1#*�8gh&��
�wh}�P$Q��SDJݫ��d�"$	�f�CM�6(���K(�"�22�
��W@%��I�p#��C��E���-�?(#�Ȟ'ٌ����.t����)��B&<Z��:�'=~��Y��.�U�3�����!�P��yc�/�o/�]�����������I�nTV�q�G>5{�������pw׎HȤ�����>gP.V@|` ��r�	�L�0����2��~K�+R��"hOj5�U<X��dZ��O�L���:n�Bm��d�'��T�{��M铿I1�6[��`sp� f�DB�%��/#N�����a!1n!E��`��ջc=�q�}�����d��\���yMu�&�eq>kX-w2��b̟��HB�I����f��ؓ�ėV�G8R��FVF{�5�{r2"�#v�
�9��mT�H
�̔B��}ҲX�C��I�o��ICn�N8�.#k��;�2>�����6��Ǳ�`�!i˅� �]��f��q�](o��G����9�e��:Ё�S��*��b�|d��E���םX������)�؋)YT.<�<Mܻ�۽�M�W	�I�h�{�X�3��wƻ9#cS�]F|��w*�������������G������ß��go=<��c���79Gu�T�iT?�';T��G���Cf/�jJ�A&�	X������KD��'�o�
2�Iˆ��    IEND�B`�PK   T��Z�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   T��Z`$} [ /   images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.png켉;��?\_ϣzR�'B�OE"b,-�����f�v��Rc�Z�P#$��R�l��3�c�Ⱦ������{����}_׹|���9���������u��;v�Ӿ
7ܱco	�{77��'���������O��X�y���[�;D>��wV;�0�Bk�D�ۡ1V^�;0�YG7g�����Yw/�D���;��І_�����D����,.����? ��?v�@ў=r���>?Ot�8���g�8�Ko��ve{��;��M��g�d��&kܖD<Йpo����k,ѧގH����@5F�G|�X��9�@�j`S.�'��[��ؿ���\�m�݇m�h��Jx۵9w���{�D�c���W��%\[����vn}����ma��������Ƿ}>�cN{��!������	�#�{��.��26��������.��qDSx�v���61H�~���/ڈ���V��|~
t�Kk���!Q츨(��?q6��k>�4�r�K)�TnG� ���*�E�Op�@�]��\�;/˘a�y3D}?��J�������%�����ٌ�<�U�Rb�pT��f�%�\��$S��J�d<�T%6��#AZ���ǻC�zs��0���?Y����z����c�*�9���ޟ(8B}�Uv��K�!���W�DzS�ڿ�¹QFn���\-�-|�&L���X^�M֫�-�d=꼒��t�?�>,�����3�ah�1 Qf��qːY�����)J�	B|U��"����;h�5횇�p���7x��-���"ǵ0�Mø��3j�3��$���6RɟVS ���Y�|䟇e��&m���>.�E�{�.�Hd�Z`����)�E��w��4	����ۦ	h��;���b(��?���3�nԛijiY�7���[�f���ʢ[�M��-o`+��]�S���ḇ)�˨4�`s��ϐ�5��i=ΩX��\��0�żӸ����Kpx��J�e�ztW�J��erC})�� ��s�>��+Ȭ�?'�a_wu޿fg��0�*�{2�as����@ۈ̥/���pK��~p-j��uۖYo*�%H�Ab$rp|�,���6�FX�0��y=�M4n�G�'�s�_�e����>���x�d�k�������f��$�D�����=��_;#�z���c��$w�����O[�&�V�
��?�ݾ��|t���A��U���à�Ϫ^&��A��uص���qX"����
+u&��SJ�V4S8(�}�")�+��i���k�<j�~-�=w����1#��5�E[�ws<7:)e�wmt�U�#g��r�1�jB�{	*C��/Z�X�����V���E�i��Z.���E�pa�L�PS��<���w��C�Q�S޹��G���)!�*u�nˁ7,�o�n���b�:u�J�����f��A��J��'.f����O�-�g��8B��$�PI�7u���;����z�>{V����K|��Zy>A5c�
/g����1�Z)6T��|�/*��,����MD�8֒��9��++�����4�`z�Mک��e}����ќ��CYI���
�Z���ŤTe0-�FY�=8����E�A�]c�uc��^�/#��F�R��kqbi7�jԯW��U1m�/̏��bh�u-m��y���W>-�2�߇	M�H7ڈ�2{N����b%�뜈�M<�S$��r�Ot��e���K2ǯ*�|�í��������'��k�������:��a1�����J�����������&�#�&W�J�(�bUOx�J<v����.��rcqC#ĉ_�E��f|��%�h0L뻸�3a}��a�k��M���<^���~(���`'���"k�	=`��5�����^�o�EjB m��h*��ɡ�{_��'x������R���f�����Zm��f�4i�U^��AT]��!���Q�UZ/E����ÁD�J+��նܰʶL�%H~�;�g��ƢGF�L?�����ť}����ōϦ��?ʱ�c�����d���^������k�i���IL��@�dh27N(��ԿaUJcmm�O��y�w=,0OL�G
��;~|�*��Kc4��M�7n��`�c\�����g���Q���I��Jg|f���v��h���)�՚���mr�)N5ڤ0�e�X}���{Xm��_�ƺ�"��%�#ǚ�a:��$m��ŗa8�$����N�B�z`���|
��q�~���A����ӻ=jić�Q}{s��6[�
o�J�$���j}�~��P�p54�!�3���A���F}�©��S��C���q��9]�OPY�v��r�Y�0�gD�0��gLm*+�`����pS�lp�����I�2�rP	~!�̕ߔE�<F	n�g��a
L�)ݽn��}����B+	e�h�s �u�L�j���n�t<,�M6S������-�2_��+@�p4�Lʾx��^����p�U���q��ҁ�}!��Ya�� �Q� ��ʪ�S�oC������������l��Okx����m����V��S}<A�mH�\���E�ֿ-j0D�:�̼Lڸxh������e�T����Zl�\7�I��n~�b77�N5i?[�SlD���6��$�pJ)�>x�ܰ6�:�v��!�	��J�"fz)QÿbJ��@��N[��niI�jZ�N`!=>��#o-(�W��\�:Β���	�9�qyӒ-t��4��v4p+��a�7/yF�0�#�j�;#�@�_2���q�B�J�Be�p��?4��j��n*�����3_����j���*�~��v���7���m5�i�!�P�V������P7����;~�M~�2=W�q6RkP��*��Z�>r�&Xryk5,�6�qJ�ϖuԎD�z�K��򥹇�+|�XP������HY_�(�X�ԭC�Λ���B0�������c��f�M,;RP����vQ儅�&Z aa���7��F�r�=�Qu;�HN����a���6��2�\��,Iq�5ăj\���n�OPa��)_Ɏ^P?���Iл�CS�� ��n��M��f�F�AJ�Q�jhȢ���1?P(i!2��"Цx
�?��iAH���I�8���5�Y ��a�|�ƽ�O�:�5@;`2,�1.&�M�hh�_��ӿ>� ="	�I�#s��ʝ����������k[���ͮ����ɗ��Y��6(�_+Ps�zuW���k�y���H�'�v�����wN�z�7���5�5����ˬ˰I@�X��&˿G�(�4�0f%��O�#�e1���
G�3�w�8fU�Y�k�g�6��M��m4��'��L����*�G�F��|]��ߘ./�t8�:oYԾ_�`uRRleŋQec|2�=��W0����<&��"��t��I�؍�6>tk�����R�|�U���񧒣a֝�,�^���>_jo�͒��7�� ` :OiI����X�C��|�_>�$��$Ptl R/��л?=�;��g��*��5�
�UN�s(��w�*Ս��ΟU@����+��*G��)���Y�x��%vUލ�X�uS�"X�#'P�O��y�_�r6JB��7x�~b+�)⑰��&�G��[K���ק
f�<�'��N��y.R,�$bΧ��ʬ�o|�:�g`�v�
s�	 �wp��e���r6�Z<�	��34U�_/��2z:rl҉�F�ޗ0IAkv�̯a?�r�b�g@����i�	�j�N�N�?M���_��I�I�KD`Re����3�z���T�����H�@���
���i��G���������z"q���Hni��}�Z�G
�,��)[�=Vi*�W�Oc�*�j.����t.�V���,�t�a��
!7S������䕘�ƨ�5d��uX���y�]Tpd��LgA���`�:xgh Wm��n���g��kȹh������QX��+�I���a�kډg�z0���n-�Xډ��xOh���b��Sa�iz���s}�������l���8X�ZX�}u�<�mpT��监�w\p�Mi>��=R��I�R0��J"U�0,+ng��IT�FG���C��ɭi�i��%���r�9��\���
Ǧ�-<Ş���C}�~����f��|#@v%cBLS�� ��[P�����;� c��=���QS��_|ɓ"��A8��6H��X�^QH��t2�nn��װ��gp�V��Ν�<qh�J� O��FIH�T�<	6�`^-(X����v��V��>�����%�;K��Ò��t7w�DPn��[��ZF�[_�8�������H�\���ݘ��0�`ב x>�[�\�⸓�i���Q@#�C4���7Pk#x����F(	�/r��X�����ɽ���D�j�| ��k �z���c�$������yiܸzE",����h�C�����b�b���D*��.�������[]��\��]ӆӊ�{V�VN��0���5k�$��Ha~��s�ﬗ�ޘϐeW���r� 9}����f��i�vn�:T��in�R[kq��	�1i�|����ˤTN�O��U{u�!{A����w:���l�դ~LҒ��\�� }�!��|\�I��Y���$/�v���ԓ'O�񰱼��kK�Z7�H�W��$���G"�0B���]"Gg�ċ]�.X�;n��6R�{��Q�۬p����G�'��f��6�:�w-��@��>�)iii`m%�^$�\��Bx���I�ŉ�xE�������N����œ�h	�+�>�uJ��D�0�@�}�����]��}ݣ�k����%�A�5j�nq�oY�\��a��Z�8EE�q��u��E͚ C�TV���Y�S�҇'�I�,V$�2[�E:M�my�D&?7T�A#���;�� ����5E&���4����,�;�4�e��̦��
0��,2�v�|���ŕ(6,
��s0�E.�Ҡ�IX_'����9:1U1"[�ն5�;���_��R���u	�F;��uQA��������b��L�'�u�'^�����J�ƀ	se��?E럼!�>���r-�5E�]��h*���!��i�#4�ҟ%������YS����J$�=���'�L�Ȯ���SƏ�
��/.M>}��\��+nll��3�,�=<~�b}u�G�Z.}��0�}" �ɹU]vʹ&�����S�FK�<4���'�]�xXZ`�T��_4��sW�b�VE�2`�b�88{	�T�AS ��Q�����,�g�䔟ck�m��e���P�
m�.��|Gn�Cٰ���TTֈX_��"��'��"JӼ0�a�{25���6�Ȩ�_�2S�k�m4V�[[$c�� �[j�)�m��q���R�,�R��D.�.%{��b"��ݵc�M��_GiJv�j3`}Ȭ�s�T���ӮMz�wԏH�O���7�R�Jt���F"M4k^���b-��5�y�fk)?��Ł
y	��x�{:��V<�r��	�5�>�o�fH�T�H��^6i|{3�,�ɞ�CV����c�T�e�8a�c��d�>��Oi�.�9��=��d�Xt8ȫ	@��a����j��H����z�.`������!�Ҙ}��U�E�1�zfY$3��Ėё�Ƀq���#�'��@��I$��d�Lk�����`R<M	6�<R*�z�7��x���jM�iv�my�?���,�nJ{��Mk��|��0{�����4@�@M�8�������[/��Q_�~-�c�ӄ���OeB<�Y)�O��ǉ%��q�L$�)7�)�hm`��Hz�
�Z��#�/�g�zc�{=�B5k`Pky�ѡ i\߉8�t<��0 6|�G����s�X���E:�$8n//��Z�A��;�� $��Q�؊t�� �Y.�bk71��K��s$��#�s�A������W0����by���vS���.P�ό��~ rK�$RJ����C��e��\:�d��W-�r� $7��R��,��(.���re4�:.N�g��g� ΍��{����!޾�99��($f�Xl?j�Z�LR�t�m5�2��gk�ɗ?g��DJ�1 �Km�ȅ��j=.
�C�$�Q���z��m�C��b�a���D���T��)9�ڇ���Aޢȩ���� �b��B�s�髬G#>��ֽb-��1_�)fw��"�G���K7�< 5݊�-��6K/A���.�*�kTK2t�������K��W��Q^�@D;�L744d�dך���� {�B�$RH]�5���Q�cw�k1wP/��}̦l��Y7��� �!���.wAaasd��~�܉���5���Z�p19܄�������ȟ���Q�xc�����Ea�A!����-��3��r:2�}:B�O�p�qz� `\�Gр���TTk�Q|�N���E�e��j��}�#x���� =s�q�R2���	��!��w�:����#�y���Km��	;�/�a e�l��J�-�6[w̖�#�.�H�Bb̫^��gO��Y�PX�o����<�dl�������igC��` ���6�Y���"��{�7dz�K�GtN�ⰦR �w�R.�-<68s+fC��Bv����Q(@��_�re����}�kG{-^#μ�����9�Ug��y��I����B�����6���.@}��R�J����&��L��T�$�Te3o?����H�c�7�ˎ�v��թ���ї��кHd�FM(�� N:���_T΁���l_~�(�8�\KW"��H���D����l{:&S��pǾY�8���xq�}�P ��i�E1Щw���,��
��O�H�D��k1��V�`JN[�ً?�t�9T B�.�4=̃u�e~�G��u��	��'�Q�F�4�h�$�5��H�q���	��%�Z��g���u	V$�o�i�ȶ������ɔm`�D�����)��Пѕm���H���t2 �q����r�N��K�������=�BI�E�"�Ͳ�ȨPU�yՠ�i$RN��	@���j��h�yS9��~�b-�x��}���Z�J�ċ�ۦ��K��/N�3M/_��,�,X��',�dh�͏�}���[�@m���\�a�Sah�����{q���ĜQ���]��+�	 ��H��E����H+P��L|d$`��keJ��P�F�s�`ˇ�-��gP��t����\���R�>d:�9U ���Y����ר�N*�������A3���� _Aw+��0�FE�Ww1�r-���)է��2�E�M�/Lrn/�I� D�~���d�"+�ާ_���Қ�w��
A+��i�wI4Bd*��e�?^01���!�B?���P���X�B�� \����#�&��4qh�������,Yy��/qQ����k#o���[l��=�c������zY@��W��=b��~��b�`�L���'���v*\��C,X��-$�!!�/����?��K�wp� �R�kj"l����-ҹ7�f�A�(�%�#���6	_^��5��f�k��ɴ��s]�	�%�_�;��Ҍ�� �1��:s!�Ν;άe&Y�e��L����$����������9'b|���+�}�)	��ሺ8T��rnn��d�
<��)�e�h��|�	��G�}c?����]���Z�<��ZZ����\)5;��\��K�%$�4�����\���i�(`� �ce���0\)�I� ����?�gs�Y/��T?��j�F+EQn�۵�Ҏ�E��ac�g�Y#��b���Zkw�_/]��*
h���S� l�Dأ�<v��Nv`Kd�_W%��y���f�d?c�\]YI� #�^	����-K�av��K�B��p��-�_������-X�/Tm	� �)`�|66�&^@�����,T����G��2/���{�����ۥ3��W������Ȋ��[$�w�#s:���Z٨(�7�P"��w�~�n���A]�BY��sB��F��럺%{�h�P���p!��!��v�����8EY��nd[�.�
�z�4`���HDa���fw��e�L�* :�L5�f/���"2�� M��H�o@��D�,=�Ӫ���\���*y+u�p�v�N���CM�q%*���v�E~��M:�"A�b�����@� Ѹ����N�� Ye���"���^
������VL��� ��`K؎�a�K%kNo-���/�����Rs�~�o�v�����3-R�}����0��#��r�i���e�i$��k8����=;<����خ��W+V��>Cd�O�>���\i%ӵ��h��Adk�b>zע���"(��5��T�u��d�f�)~}F4C�#��)"���FsY+$Ҽ˩Э����Ъ�����e5��A�U��'�u�VCj�8��$���[99h U�J�A�,3��0���Z�M��m9�\K�L�]e ��]M7a�?��(J�c<`w�s��T+O�s�^XMi��g��?�S���-��~du��V�$�@�[�9 B�������^��%���H΄���<o��֒,+���~���J�L�U�ݻT,��+���؞��G*����Yv�]ߡ��ɲ�~�tځ���[s��5�j�	73�{�-i�(���P>�[�KMS_K?ӴWѥ�k��矠!��I�Ǳ�7J��8me:���pv
A!��]��2�	M--��C�nB�3K�>/Sai@��=מB��J��I$I�]����9�I�6qi�a��m\�_y]X*yrxC�?�T�$0ӄ��O%m���fAC����G�@Vo�a��gO6�e�Т7�8S)j�|��0��,>�~ z�c��r��k���ɰG�@UHA�b�=���OF�2��=��H7&�Z�"2�$�q�]� �G@0MJ7���]<~�7�teF��P��d.C�Lߘd������+��L����w%X��`�tg���}����L� �n��y��
�
�5���WVn�/����tӗ0O6S�O��9r���w�O���u����A~�2X�j�Gi��Z�(o��7_���D�����w��H��(�$���`��	�6U%�lR��[��T�;�k��-P盇!S��Hm��Y�W�1k�?�M��n�
ǁ}9�6�q)���+MM��2�;õ�y:
v��7� _q�k�'}V�c��,�kV:���]�]�P�_ld��ڽ�5�*6\�d�A�ö�(�"LL��9�F���-�Λ�(�f4�F`�e��^�Q:v/��trm�Y��`�	ɓ���d?���x��S���ט874	�5�]Q�i	��N�A-�R��*����t1a�7]Ry���yo��b�V����Q�1m���i��"B��A��ݾg�u�Ud��	�����pDc���!@�Hn^��_$��<��&��p"��)��(�����5VGZ�I�����A
}gT'����F��11��ͧk�m�N�׫F��4��I`
(&�0?X�Y��`-F�7���?3��n��(���< %�X�Qp�6���mM
܎�D�c�(lCo�}&���9c�ȍĆ�0�Ȩ�='%�eO�{����wf�z��y���î�j�F��&o��x�Z�zMP�6��'��[�w�t�(�BB@2��:�A0�v>;4)�8�H�I�8K�Ȉ�Ol�Ě���:��P�+��Z;$r�K�y��{����8l�6z���cn�~�{5+��`��'`���yo�	\��;\ó�"|��M���sd\�%d�;��~=�L{6eᰋ�x�4��,�����k�DH"�<iR�!�7Nb��;�x�5�s����a��Du��Y�Y&�1d���v����1ZE^��6�;���*��7�}�)v� �?�K1�yw��8gr������n��b_�֠���V��!�{1�ʊ��X��M~0�&˞� �S�;^��t
:O�{	�c�nƍå�y��/qLm< �� D��ôgh;m���V�����g����Z�"���v�ç�eN��D�n�8/�T�/��]K�/���x*� q�C��&:")����!�M�@y}?������G�ث{]�c���H�l�����ɵ������ɈL�)�t�C�+c���.5j��|z\)`���OC������c���+��C��?J�)ʌ�@���]�3�UΓ���o/�O���%���l�E�Ѷp)�,�ɜ��|�_W���'cX�YD�;eG~��Ću�0����0YѺK�s����Ǖ��MesU�QzD\�B��o����	}��1`�;���ՀCBҬw�����U(�ΐڣ�����?��Wǩ�Wkf�[<���C""��@���VN���h�����= ID`x��W�6�8c��{��Բ�;�7�=����LV��&y9��҉
D��YUl�����h~f�jg���~�sU�n�5� "{�a$67Ț�����uU ���7�E��;o'�̹����_}x������e�D�_2G��S���y�÷�[��>����`��n����rN��
w9C�}��9(vH�t�,��V�>NPX*Y� 	��W����XZ=t8�*\=���y�4�G�fu���e� ���5*�Z�Y�tl#\��5d�+Q��/����V��l�`ĸ�{�7lt]I��RU�f~�nտ<��0!Q��<��x�NF��� �ͱW����]�=��k5-������;����'��|L�(�m��p��j�^'������/���Z5Q Y�����=��1�/ꞃ�����{/���s�Ĭ���VDs-������{OZ� �T �vV���2��o�C���6.jj����%�t������XJ)�	�q����?�4����2�$iv�x���X�FxxlN|;M����������F2f�� \E�A���j�-�DI-�^�B��A�����	h*�Y�lx��A��	]�d7����g|�8Ju��rƩ{K"f[���TF���'	�HƓ Ti"�D �,�##���,|���ԛoO����و7-D��&�U���l`�'tt�y��\��A�*�$��]{5�� ���5h��	�"u����"?[��: !D���3�����@�Y)JhU2Su��� J"YHH�g�뷙^��Ei�U\u�F��B�>��ް��F��������j�1P�ғ�ّ�@/ʾ�g�b��>���bN<-
�����e;���S��Mi�,P��8�ͧ��n��ڮ��"Z�IxC�2.;���F��s�Sp�ǹ�i�k��'���y	�3��X�C���W�
���h��3��g��B���s��'슨Eٝ��g�W�T��ˉ"��~���L�,l		���#Z��uIS�Ep�O�������WeP��֤�����F�C�ܬՙ�]*�����e;�껡|G��w�%�S�w�Ş��pǏ��*�1�S�U;���(�����*HT�W5��+h��:�/u��D �M�[���T.A������pϭ�/n��{0(i+zx�>�[�������$��u3�}�q�XT�k4��M}�(�������4{GJ�X���a~o�n�ĎE�3�-�8Ne�j�*�_mg����>p���>(��L3|x-��f`����p!p��+'���N��x�{�M�$�=�~JC��^��4x�l'�/Ϧ^�eԎ���+(1��YQsγ�9�d 9v�*Ψ�A�n�P���8!�1���H����o�P{"�3����<э����޹�7-
a�^����\�;��DJ����E�B�G����;O
��w��FJ,,�~pdR�x�=O�����[� A�T�M�NlB�4e<�S���k�y0�#��+=3F ��)}���Ϛ�a)sNm_�lڑ`�Z�x�-`�/9� �[��l"׫���d��L�Լ��L�U�#�^��5��L��J9��
h'�iij�Ĺݣ$���q��tT���hJ�͡�n�.��ەq�5�Du���Qʭ����ak)�b�
5�y������*�5ۿ�����$Q�c0�P�M���^��.9�r^�����h7DLL,�����=�U�
E)?�i(!g�+p�UF:�oZ���Zp	����7�JˍRhk,T2��D	�mkk� ��oy���������E�c}���aC�d�&���aZ�q1%Эzgؗ���.+�ܩޙ2�{|�����}+Ľ�� Ǯz��q�;`��������zRB%���R�ͯ�r�=���9R�- �^a�o~�j��)͠E&F�/�f>�%�> N܅�_c4��B�"�cajg����-��ph�FʜR�_8�֋��+�:���ޝ�+��FY���qnY|�����=�V�)���;ĳ��+�����_�H/;�,	�￧4����ؿ���D�T�+n�=�W+���F
����=?�d�S<ـ�Fuv�"������Hq@�>g&��^o�Z&�/?���f�%'�Uٱ�e7TԚx?Kb;�+,�j'
����p=��eN�d<�w �S�E���$�Tn��6���J� {R.��Cvˢ�T��=��JXJ�J)u�u*����؛7@ϔ���LKB�J4�Ji?�.'���<`��-�S:j�Q��;NL�ƹ	W��s��WM)eyEC���3��W#y�t�cz�*x��6߃=��Cc�MD���5W�?���8[J�*�@K�˾���0C��Vh�x^��[�s�����p�	"��D�I���K�Q!�s��P6o�w[����3��)./�ͩI�~��cH[ʕ+V	R�>�xjݩ͊��
���dq������;����3t����d���v���8U�ک>�/���`����,�~�?�}������P�	 e$6lo�o	��io��K��H* e&d8R��f#�l�׺d5yn֙�߿��j����U'
���DW6,����SKU�m�'�4��U�`jF{�٬�#ǮJŶZ2KT�(A���r_��KB������o<������V�y$�-�FE@�.<�-��撐���r�Ox��aWZ��&��Gt��L���!U{��t�h����P p��ȡp���_S���#�<��X��e�ƩC�Cf���N8���ܕ3�y����o����a(<<�`5�1������j��>�A��j.�[U?�Ҫ���	��[�[���
��`4
���$�Vl�[4��j�v�ߊ����7m	�D�v�(K	�̻��l�-m��y��R��4)��)�Ӫ4��]�~FW��[7�1��N�8V/�=���Fr���EwP0L�R��R���t?����?�9�Հ��xR�D9�;6"��d̼Z�O�F�&t��q�|�ʵ����Q����`�y�d�ܨ<�+�=�պ����f����.��~ԭ�(4�������z0^�>C�Y�pB��� �����!έ�H�1�{/��h�2+�WX��*
'߃��P���_��}C�Ȉe	�爝 K�ɕ��j�H��!�����/w��l=�˸��&	X��
�f�>�>��-�Ů���حP������|�G[�� ��t�D����է�aw�} E/��)o�X�н���p�9$�%|��䩃BH&�s�#��D�=\�
�5�6=o����Ha��!H{�m���'T4�6� �.�DJ�qq����(w��N��Ib!�H}���W��[��� ���e �}���[S;�b!`���?{t�PbXFa��w�2䡅~-�52�v�l���������A]�ȳ���6l���� J��yL�90��5B0G˽v��DGGFbOaOb�+d������� D��ֽwd|��n�����`2���e��8�!�����T\N<��BZRxg�q��x>K�)_�z�P��ȼ��΋Ld��S���q�w���� ��~������U7f�Ǆ��X�{��Ndz�*|0���{�S�͕�%��+�`l�_���<ȆF͝��i���?c~?�pgaz׵4�(�ek����p(�jআ�.3��X��z&��Y1�W��^�|�'G�K��u��T�#
��.��7�8�p�hY�r��Ӟ�l��kY���}�19�o��K�F���OKK9$�I�H�ir�F�Q�Bt9����B/pl3;r���P�ذ�i:�sh��,u4Km�W5�f2���	a�ك��6MF���p,�d4�D����b�N �7$��\I��AK	͡s���%�z��@�6R�Y�'\� �ۡ�� ��Nף�F�,S�ᇺ��H%�t�n&6�������� E�~U��k?���lt0Uw��O�A�b؉p��Z��`���� ���|c����H�[/4�g<%-$��Z��۽��� ��J��0q�\�}2��s&Y�J�����9;M�{.�Dw��8)��$���+�peҭx�UXFȕV3�����f���䡝zc��|���RqP0H����X�~o'F��G|��]���nn��jľ,9!A�������o�}�i1�,dc?�B�="�7��\��H�~�#��d�A	���~�J˝�͉7Y�/��98W0�����c_y����~�{�Me�s)F�Nw|�=+��u͉��>��m��(^IN�=��U��D��F07%�V&Z?{,�ަ�"�{�}¡Ё�b��Oh2��p���j�C���m��RwښIz1�D�f��P�OB����ٜ/���s8����P^����l^ZZ����E)O]#x���`%�ñU&�+�o�uL�i�/�&5�VTS�8�D3#�L,�	Y��b@f����w�]��#I���sO�d!�����C���/��ۦ�V������~�l��gŇge�cā�{��tV<Y�V�S�w��w���LsPN#Efi���TN�]ܹL��v��f�kkKU}*mF�0��U��f�7&Ai���B%���yy#�K_��t�Nu����H��KWV�M�����	�ǭ?�$�6��_�et�A(!9���-"���ʟm;�vK��<1;胵c����!_:��
3R�q\a���d\*_�y�����M��s1�p�&��)�y�@�����`��� � }�V�ʒ��+�~,�A	�����/U9?A���n�_�)�v[���#��HB�^�Ë��_`�"��/�������2�8X��)���֑H��|O�:1�qLD��=��*��L�y����#I�&���X�=0o�J��/;R1s�Nns�fݰtc>z{� g�y�ʌ�3if�ʵi����61z�.����RM�rvN�?=��v0�:�
R�򝟨��T�LJЧ�-�a7�Z���LѨ�D4;�U14�bo�r��"���J�ce4Ɉy�P(~Q�a^�5�i�Ŕ�V<�0��ڸE�� �	�j����3�'�]�_���'��ڜYbh�ᬚ�L�lÏ���"�{)===6F�S�-p+49��>Z� �c�"�\���ߐ̜ۥ^���{��H
[þ��,�}�x��Wf\�n�X1�%�jr\�^ ��G�U
�MwG�Ś�e���Zd���t���Y��G�b�*�=��YqZ5qPkOf�v֮������:z#�{�(i�9at�E7Z%������e",�P����(i����V Q=G vo�
7�+1
�~y��U�Q|M#a�=�l�H�b�ᖞb�ɵN������b�^��Z���eO�wn���T]��#�1��%�@m�C��ʄ ��Ő�U`Im�yۣ�wj���=F��`��� W���\�.��/x8��%nt&ʪ�B�}�R���<*+�o�']I�PB�$���o������lH	����%9��.td"'b���I����ӏ�1�6-�{��9�t��`���wU����@\k�����a�ߘ����}�R��j�_�n5�߻m4=����	�
�w*hg���V��+��^��{\��\�G��lI	:�ؒI w�U�@lXf�3i�[LI�����\5�������a�}���M�/�9��R7V�QV	��$s?μۈ����!��lW���G�3�{�7����×��z�����X~��;��!3V�9�e�p����xL&��ʘ��t2&��ovt���L�Oi�2�c�*� 9����D�9ʈ&F����3U����4?pyT4
`*Ԏ>���]^i��a3�躂�������$�i�eؼ��5� 0�����sS�Y��,G����%Q��mLg�����ͽZߒHQ5�`���ȕ,K�����1F�&	V4`$2��k�}b>�c�+(E?'<�w���6�H�C&u �,P.�SheFDTT����  eS���Q�ۉKk�e�-�}���H(���v�8g��s��̲Y)�L1���~�Z?sR��*�����a (��uۓ�'}R�����OV ˞�]N��;o�/�U�7�V$ �"�I	b�1r�o��1Y�A��:0c��n�5*�hy�4���X�V1�⩵��)�iHd�Q�^�I�ߓ���̦p+���#�ޗ��Gs�#i�x�q�Y�N�r��Y�JP�vCj/��S�Kѵ� �v�8��:�x��t*팊Y�NL��mtT����wT�GN����X�o�J*'��B��R�o��_@t�Z�y�Z-��ksy�6+�G�����4ۗg(=P4W �+�W��/���BG��[viX�r	b�伿h�R?�o�T�'�rB6J�-
�@�$�:}1.��;n�)�L��sC��O���c��~��2�zKׁLw���W��ݶS�<�`���6'׊I$�b���Z����	�b�~�X��)-U^��/�xh��� �۔���"Z��=+|Yȹ���-4L^��*9Mm��6��{���W�� R٦��s�1Ȕ�P���y%F���#���R_�{���Wϼ��87#���G2��S�TDl������X|��E0Mt��}j4�n�����1��6��&�ؤ�<�g���D��矷�c�$�$�Y�Ԥ�+��Bt��)����;����cG0��_�'G")�A��%��"&��_�fv�+X}���ab�:[ؠx�D�&C%/g�dmvfr#�7�i���Ubl�*�Ք��Q�63h��O@i���sr� ?`� -��<d�٪:QvI�L1i����X�]���c�;��o��d	)�i����(O$�>n��({�����ғf�@��+G,��ʧb[o^���g/VD� �W��v�=RAW*Wp�C_��I���TU9�Ҫ���۫���;�}TK�m=�,�BSl��E�"1�"�R�	�iVBƭ�-�%��\�G:@2����q�nx�^�cG�b�\�&l��	��8��r�7;(M?�b�E�v������9�07��V1�J���uoPF�bo$Rj���J�k> �O2ި��0��ĝ����S�H��Y�Lt]���z�pmX `��D���$	�O�(	� ��m~�-jέ9��½�w))��?萇���_��h�{@�j�?�wTS[�.�9�=��5
*D@�[(
"(M��H'���(��
H	(H�^Gz�R�B	=���������q��~�x�=����lϜ{g��L�n�٘�@�/��"�O`m1O�f;Ύ���r�u������b��⽨�g����sV�]tH����_��s�
�8�wY�Q3���,�� 'n�� �'�9,Z�A-��I�
¤F-DےS�����1�}u�s��~���^Ǳ�[�����e�=�F�~y4g��[��۳@ً�>2x��Ϥ��Ҋ���7oR�,��]M�	}��Φ �|�FOR� g��U�ünۣ�����qZsk��h�Ѧ�i��X��-���%��W�1g߸��-�/p�����$����}J��8�G�.������gd�(<A���Z��As�d�X*��*`�1���[�.ݞ �B��#%nv�gά�uH�A�+3��P�k�����O'��&_���A��Km��k#�,0K@wR&�[@6�T�M5�`3�UϽ��D�/���J{HB�4�����Q��n
X K�t`^�k��5�@�t��z0&WU� ��*~�z��η��-{�H��vi%�T����A� Kp�t��8`I�:�f,L��%�3��#~z����aР�����7Dɞ��1��5�>��F�L��=�
h�4~{�·�۝�\e��]^$2��\� o��4	�k�Q �""Co\�2_F3���p97�z���*����C����/��*s��6�B� 1��lړm��5�l�0��(�>�Zl�'�韼��4��L����?���7���Z�1hQ��>����V�0(>�GK0�09������XuE)s� Pf�*�]Qq��d��B3�/:b555s@��1ϳn��8�r��3kޖ�b�20;��9N;��zވ����ϓ�+,%V����Ҋz�,�>��L���B u�dd�D�b��V���`���":�\u���M�� ���|e��b�/�]��$,�6j32tӠ����w�whvM7 ��Қ��R�K�� ���~���~��F
Itն������U���X���s�8v&b���A�H�#Yz���{Z�}�Wu�ں��U�����ҧ����)T�@2(w(,=�7��������n�	�����n� ���#p����Z�L򇒌�n�����f��E��@!&y����DZ�~�/�[ �$� �#ޒ\�;��f+'�35�K�K���`�gN�^�7��n�|B�UM o�ǩ�{E֮��a�c8�����\�`���ӹ��G�֓�������Ѝ�������7�
�V�Bu��7*4���p�hOТɫ �Y6��R����
�'�����I^dg��(C��n��~; �q��H04$D����m��
�22������i����p	��nRgg�+���휢���jv�j�k���z�Y���+����v��[�|�C!�
���Pɚ&S�i���nR׎�����Vf�2���9hw�I�m�#�=���Ô3㪐h]
�4����t. ���`�Qf$���#�`��H���Q�[r�T
9��f1�����/˰�V�r5��>��F/j�6�b1��KQ��E�'��,��95yݺ
:��n�&4�E�8��)u@W^>&�V�H�8�/��K��H�O��+ܕ@���)�[ W��k0n�kǗ�Sv~SWW�i	��uie��{=H�XX���:�_�Q�4��mCG��K�3����L24PK�Ȑ��F���kY�"Bc% ?h��.?��$� !''x*�E�x�q��e!p��&X��7���(�1���R�H��h��eZb��&�u�k���������7��US�K^ML���p5�\ݒ�U�>����S9��A�����3���a�~cZR�Ǐ *w��r����[k�m7F�pC���@����^t�W�hT?{a0�Ǧ�K�KTO[u�qp��m"�: |}@R��Ww&��.&�Fy�P2�)h�͍�"\,������#���PE��
���9��[�<�[�3�x8���3�$����j�Z�-|��w�a�k&˷��jU��hU���{h�<��	-�����$E�!�E���9������n�W���cj�"���$�o���`�c���+�'�*�,q�n���ļ�b��ǧ;d��[�)�+��Y��$G��e�r�����}T� Ց�%�ٱ�.�Pӎ�ã<�f�Vn'�Ww���W�f6]��R�4G�[6~҇�s��vôS�p�
���k�O�V�*~�I�����d�����&�#�.	�6ם*�j� ����Ama�H�eR:�R׋����<��F��
�:�?O����P�AË�T���+5c���-J`��+BI�dS�����Z��<^\8Y��٣��TMM��Tm�	�	;�d��Ŝ£��f�b���@�KPQ����$#u�\mӓ�S�<5#*T�U3��S����%	~>R�)�v����"�����e�x�
i����X��H��v�:i~�@��95j���?�f'����V��S�?̩�7�U���RA��&��El��P�{Y?َ�/?��ѭ�v��j?αRe"�2Q�f?e��(��~�A�U*��l���]��Z�VX������� �����RO�z|h���l����O����Y��N�IkG}ۓ��d�t@B�4g��tm*\�u=��O=������*�����z|CP�e����A�R����T�� ����.�kƹV�hΰ�l�,oY������Й9"��W=*@�z���9X�s*���X�)�-df�����'�/8��T]T��|��|�C�!BǏ���h�����<Ԡ>��u�\l���yúQfX�T�VT�\_� �T!C�8�c�n���>":���S1ڭA��g�����h�.#�1�H�n`�1,�g}��E{��DL������9q� ��
�s0�Q�����tY�\`T�a������OoS�Z�+zJr6xxG']���t��g�l{����UH�+L�Z������I�*.�j�V~���
��R{:��~~���#~�0�,/U
�w��-1��Q����^F���⦵�c�Z��û���=�{�6�� I/&M�;r�1���
�9�FU�&a�<;rgbD�`�1
I��}	d5è���I	��$���}� �����[�f"�|���O݈�n>��DvP��((#�1)��G�����.:�'���-X��,�h�b?�$>����:B���h����8���VE�ߡ2�����Px�45�W#�<��¢�e�6�p�PO&�8� ���;�^`��l{�jFur�P+!@����c�d�=�P����Z�3,}��h�:ի�in���Ɲъ�	��?9�JL���wjO��iL1����O8?��vrN:�9T>4�A�v`�{�^�
��%G�^�ގdo}�\��~c$�]�:���k�j:��tY?��-�zδE���i���s�j��UN�$R�U�A�h�^�0��K���[yB�.K�g0R�lfZb����}�۫7Y����+������L^�d�U�)�E>�\�ں�1r�vB�*��HeJR9�
��/� ���P�.�J[�Ti��j����0	����UV>��m?P�|�����5e���������j�(	+;B��� �S�=i�::_
��H%Q�5,6a�	�Q���ѝ���%ahȥ{;ԩ��An�c�����E	����Y�s�Y�%�Ws%�yb��ˏP�㫏W�OX��/ϗZ�焮�-��.52�ϻ�i�'��w{��-���qH]=�k���Po�G�k�l��'�Sb��\����%�& I��"���,��^�nJSY���'��c��DdA�(�,"ɐ��"��^��C7h��zW45}֍9M��Л����IG���'l��d�u�����4��]C�R�Ϣ����� ���A��$���t"�-S;����,g�SJ)�::}�4���S���m�����B6W�4��K�ȷVb���]�T��9� z1!iE�Mܼ�'��1hj�3I��j��?7�.�F���U*%>�X2 |d+	�g^��]O��O��n���s�ǓHǝی��Ʈ�R�uh�g�I	��3.?I���B�V?'���'����&&s��+d;��kx�9��w����e.�='߂�hC���+����ь�M|���)d
h�2�����/u6_詹4xI-�	k�m�s�]�_���֙T��]��g;�xs ��ޣ�����)��$ �̈XC�3V���.K}Olt{'c����\Nu}�%+�n0#f�?��T϶�̮&�6�s����N�n��,c'�/?���j�D�Y�	�ʯS�����Sོ��"W;��C]a��r)���3T�v��Lk#ߓaO�.�4��tk�u5���(Kܲ]��Qû�e,��Q�q	��N���v��nn����d9�D��\X"�v��Gt�~����X+0�>��mѴ}���Qƃ�.�]��8��'����ﱖy~��.�԰m��ڇb��P��W�9Ƭw�^[5u����SexhZ���Y�Rpj���W��Y|�%�\��(���i���.�����O;�c�s4'��߭ �W3����E(k��a#A�	�D��c޻�K�|A��Z���l�U5:�м�����F���]�f��sgk]m�Cx�H�A�M�������\�b�Y7��D/��k�����~%���z�|M���&��ߩ�Pɪ�����mC49VH�2�$P�HX� ?��=cɯ�q;��koT�<�$u���*�8����J=�؍��,p����)M4�5�~��9�h��C�"9;.,�J�:�[n,	Ȫ�%F"DO�?QcrGN������n(�'�{͓h?}%⁪[F2��y�����$a��sI$~�V[�����������[I�y��E��/M& ШR @hUBB���V�U��_�,ñ��Y}[|`#u��lI!�xϤꣾD����ѵ�1N��B߁�`7�*0b�?)��Q�?���V*Ur��o;������&��6�nx�W������~%���q�r�g����}`$�L}��^|������s��E��}�T5؞��䒗��i٣1bAەx}�E�;����c�B��I!��jHMBI	�q�$�p�݉=>�.G��O
|���9�0���wB�� |��IVRn��1q��O���(��GzSS�ߑ��\Y	'��1e��G��T�Y<3�,�E±g�����S�U�.�����VQ��?�>3=����2�O�I�\��27z/�����퇰��	�I����@tl�}�f�<Y(�$��H���C}���М'bߋ�w���p�l��H|=i!��B�O��JlFT��
���!}a��w^v,�
�����adݷJa���uy��_��yw��3��H���׮�Ɨ�,tܥ���������8��ɲ?]�SD�b��O����'����_���O�	���>���K21雔��[�G L})�_�h�C�K7-#FQ�Bydl����ձI��p���X9r�^A!i�>�&l�󱦻ڇ���[�Kuaj ������\Q�Ln�˱�uhU]��RՀ~ f���c�CjK-L$�б��L������Mu����r�y��8O�� ���0���ϭEWpy�Q�V�p�bg�o��/B��,�<��U���z���L>���P%��/<�`a(���ᾅ��L�p�*Oĸ� �ơkR����O���&Y�W���䩀P��ꌹvP�q]�BR���AgJ7����#�4�'����-	;�0ə��)z��9��f���	9��Y3�k�KmZ���jRީZ��.7���gXQ�a����u1R}}b�"�KY�U)>�_�X�u�b�����KI���d��M��uRO�Їf[khXu� ����">�%6�Ay�$���p��`�t4^������+���]kd�n�x�%6���&�?�����UT R<l�jEz��^���x߷��by�j���O$��|���ގ�	���26e��9���rΑA�_RGC�4��۽/h�U�~��E4N��$�À~�/`\���� �W�ǽ��TE~yPƯ�2��]@������W���
�����(��W]���(�����rH�����ĐT��f�����R�=|.Y��e�,�4��O���8�8)t�Ƈ����+Z[4����ꨁ?>�D$>� Ѡ^��Rkvw�q�i;_
������W^��ii	g���O,V�=��R���Nrs?y355�'��א�]^���%��%4i7W��KUX�g�dgn2ִ��x93W�
K��(��LDڟ�<�V��2�Q�
�A4j�-a�����ȗ*F]�0匈�AnJ}Ή�֔h�[���b�9io rF$�U���yRO����Zݛ	����p���mHn�,�~ms_Q�?���5��ncoxwC����4�Js^�>S���E�l��#�d1L���Uk.U䬭�Ʋ�V�Q������D�����ƿ s�	Y�hzY����
�C��;�I�0Ǔ�g��
�ދ�������_lJoj����+��5{zd���}���w�P�u��/���	�X6r��2���wW&��"z��CS��matt�� _zx<%R"L۴�nҟ/��`�K����~]��y�V�H�v��䮏�q���@����=>vQ1�J�b��"$�6���#9�N�*���9)�IP�1O���	0�wrs��/k�cs��;�]��,V�;;Re�Ml| }(o�oh�2� C��k1�c�`���K��wk5�[��^�4>j�][6��8��t:G�io�f�'�C�Ѽm��t�������3�c͡�𕀋����6ѱ:��W9n`k�p��7�HA�6*ʾw���J��4^�[@re1�������)/�U�~6��s�d�^C.X?�S� 'Yu6�{��=���^ޕ ��u�Nz��b�Pᇔ����^�{��9�����Ǿ���������kJX_$�P�����0�^[�f�pQP9�3*ok���0��FZ�N[����]�C��z����9A:�*��t��>�B!ij���x����<�N��ǎ��l>o�1��\t�����6
��?�����
?Œ:�o���[W^����װ��+'��F�%N^�Zu��k���:����P�6�P��=���K9���
^gx�[V\ҟW��^x�Ԛ�%j�;'���C���q��.����1K�*��o�'8����Ú�>�5)>��$�;��ܧ;3<+����V�2�سp.6�I���w��r;*��DL�(����]��2yz�@:�7ɍ"!���u��U7'�t]fbr�=K���!r[䑳˃��w�>�fhA���j+S�Ǒ�
Φ'[����<�Q�(�<Zc/A� ��8=��Jo�y��J�od�W��%z]ɽ8��3*�w�g͝�F;�2�d����-���t̧]�	:4�QΡ���;��R�&�
e�`��4g(�W�{�&�n�(���F+$&[�m�S�|YA*M�=f���U�D{$wN�*Q��O�Jw�+��o�N��6t	��s�N*M]�o��㩶���#���q��▬z�א�ɻ���Ճɘ>Ҳju�.a�v��me,�=��CD�\���kd�8F,�"�LQ���B4}��6�$���qV.yw��p$���T*�S���䗍mA\�{�`��gP�v��P�L��*q1cl�P����yF��-ʊZ+�sn�+����(5���<Q7��_�H+��C�2*>k�R�Vn�%�r�5U�L��W��ԦV=I_��y��|B*���l���"��Ҡ�B���
��J�>狹i���O��TGcG�v�a�on%j����z1fk���@+���Ɖe�@����������>�&����D�^k��x�3�SIPH�n���NU%��BjОd�p��\`�2�`UP.�u���jP{�]S�N!ӂ�\".N!��Y n��V����=���D$Y�>B�}�>�J3��'��/T�]�KP� M�-0��J�$��<?�K����j!��E���ڞ��^ǭ޻������A�5q����i}���^ͬ�F�|c�f�ω'��Z��w"�Y���:3��h�4m�H.)�R39Y��u�T*Te��ګ�P���T5����<�X �̃Z��$JИ�E#�㳫�����	/�x��-W
�KCJ������{�e�a�����n���y�d���<p���z����f�� �:́0������ �}�D��`���F�PԮ��L>��0D8a�\�y<g��e�h�f��?��T�%|�8�2���5�y�_�VtiB�v�r?6ʀÔ�ѿ��d\��jy���ڟ���ȭ�P6�F+�١>��.�ݥ��;V��%��������
��AC[��I�@[����¶Y�ĳ���t���:�����&]��H�T$��9+(�|muD��Df]�V�]�K����P��>d��0�[֗=�|��ZXi�P:�܊0@8�CM5�=�휎<n�A�x"�:=PT����1��ܪ��	/DfI!
UY;�K��yy��5��W�m��1�3ߑ9N���?�(">��LɫUiA���Q]p*�(T׫�S+ז'������(?���w��K� U�h~�e�.N�6�C�9��K�P���T���p�V��k���vC�|�xC-���;��׳th��K���$^�y8-U�YW��L+o�l;��.�ڪ��J ���o4N%�����7@,����q��~��H��G�s���8Q{����ar��ҭ�ϓ
{Ctdܯ�D&{
���#��/k]p����	;�r�7�@' L_T�Os*#	��K����:���4���.��=�Ჲ���J��k����Wx�e3_8���W�;Aז���m7��@�/�%} ��qA
"��	d��_��d ��m�kc��/�yyｯݬ���f{�#4��´����|_��b�Ԅ���썄6q�&��O�T_*<�{:��I�]��]�yk�
o���Q��8�=t璠��S�ow��w��w�n��~\���!��O]�#*��hq-���8�D�C�G�q|�Og6����v�����@�{�;R�x�lŃ�/L�v"d��S�.<�y���g6f�^1���;�E~A�~�%�s!�#U6^��'�˲����U:)M�u��La�fY���k,vU���:n�5�U�����H!����M6�{A�.j���ƫh�g~F��&�k�	؁����)���˽/���b������o�Y�̚����˫hm��������.9دeIn.�F��oьY�r�Q���T���K�3�2�x�-�oJ�O��)�)h(#MCK�+6j�y��O��h�0�뭱T�w~�%�Ծl_�j��8���'���a��U40�!��ܢ��5�����j��EQn^m��Ŏ�bi��`K��CCǥ[��l���)9oCt��L�L�!�v�4kxa�4ܻ����X1�(�YU<����O�
�^�s�C(JkGjX8��d� �[�)�5jiU����ߓ;�_�7�۰1	��(M�76�4mё_$u\Χ�Q�#�&��"�#��_�LY�_	x�������\+�OϿ,����G=�l�բ���@{��+��c�O t�b���涮S� [��K�L�e��|f��{b�q��$�eڀ,���p��n`���`�
�]�
`t�fփfE��!ǋ���7��ц���:t$��~�;�F��-CMSծ��X������ǊuT�_�c^��I�FXu��b}!ڽI����Yk�VFUD�Fl@��Mٰ���k����)�S��6�����>��ᯜe��i�b*�CV�/]��+Jpu�%م.�ڦ��K�Ӊa�7�M1 �L��g &
0��9�-+��S+��Q�&J��㗍����ߧ%�~m��*@�/D�a�z���"�y\�X2�Ok�fQ��7�jB4�[�s�ۚ2��k�r,��t�usJ>�34b^VuLu-�*y�c��W<tyʪ0d8�`�٫��Ĝ�2�;��{z!n��P���c��Ȩ�o}�]{䊚�h $s|`M�R��i+M�����3}���o�%���=�v�M�iŕ\�SV�>?ZL�oY`D-����k9n뙈zG�k�V4���K>ܫ:`�]����5_��=hC��s�Z�Ɣ�y��ŔX�e�Fs�	pV��0�w=�ۥ�@��Y�SE��a�I�&�i!ǜ����n]KXy>\s�ch2�Ϯ�ޡk�1WL.��5�λ����<@�uE�0�Xpۉ����Fv(,P-�@��".\�����\��ܼ��%�<�X1�W*>�C���f�'�n�߽����<P�{ ��[]&
ľ4���A�[y�XP�Lz��XJ�����fu��2�M(ׅ5�A�8J=��n��{-55����[[�����z�J��Jj5�D��+���P�dQ������h�5����"�a-	6+�"�UHTm���Y�y��u�FS����v��<�b9��=v�ѡ=љv&b�q^�I&MZ�0_ւи���XT��e{��5��aA��>� )͸����V��v��go�jD,�� pH1Z�L3�Y׼l�<@Jս.��`z�*�hJ�I�������|��E�I����`�$���w��ڡ��\<��6���}�غ���sA�'$���!=���2o�|	���95��һ!ȕёb�}��Ux!�f�e#J�}`
�O��+��"�z�N���N�θ^cb�)�|�E����Um٨�[B�"���-��))_����f_�3�漄��w�n�c�,�3�vN�x�(�-Ξ�9�"0��e����F���;7��?F�L1� �6����X�YhO K�Z3!�..LK9���g��A���[Q���|��\�#��,w�H����ۿ��ލ����m�1�}y�mÛ$&��q�q�:��8	Hҹ�j���F#T��⥜r���ue_i���8v+�vt��S��8=�U}#Pu�u0^Г��_-�=��*밼�����N�f���Р].\Oy.h ��s�P�h��W�����Eg7O!�}�>
sk��pZ��#ﵬvg�o�����htg�[�G[�|M8j�9��gby��A��������Қ�Fc8t��3/��U�(��/�X�U�5+�R�ǃ6�>�����N��ɫ�斖� �&ే&��4��@�[4���X�-r��+������Bl4c����	�X(�r|kmߴ��pZ�ޣ�zg:h7��\gem���&GGϜ��v��?9HH�n1]�dV�*�o� � @@���+�Wt9�^L[U�KB3�u�Gvyh��-4Ꮚd�T������Լ;[W�fX�(�ƣ���F�k�z5B�TFUFO"j��#�e���-��`����Y�o|]ׇ@��{����ަ�Ym��
cNIM� p�q{�ln����v�85el�RP��$ �<���u�!d�$���HO��44��o���U��+^����Z֟��;;��ywi&[��m�Kx��G��8��ӗ���R�X�9Yd8�����g竑OX%�D�Fɉ�+�.�T%pY�i�;�4�CT�U4�$|������v琔���J'���ͭ�7?�fЭ#U�x/��-Z�X�Xi$�����v��֭�Ĳ�'�"2J2,Hs��hT��|҅FJNMM�:a}��Q���� �[\\�1Z^�d���ǘ`1�! �o����'���y�I�k��j�f(�Ccs����ZG�J{�YE"i�����%B�9Y��0O�]��J�>mh���y�����`O��4��Y#��xs癱���v�C���9Rr��v:s�Wʶz�z8�N�DI��y���snD��+x!kr��&�Jkh>1���tΜ��7ă��E����өa$>���m8��f!n�����t�Rn;��@���iGb�9K�ݡ�Ϳ�%��l5l�mN
�+/^�F��rZ������4�#��}E'� ��\��&S'��n�y��lN��Z=?�����cY��X��� �IAN=	EW)�G %�BkP����P0�ۤ�u������'@�+�v�lg��*c��F{h�p�{��u/_r�a<ދ)'�X@�I�����U�����]�n�2򜎔�+{W({�N,�Dj����O���B�����H�qJ�4耓�:<@S���f����/^\���Hx �e��ܱ�'-��Íh��H�M����[Z�F�2�۾`�]f.8��m&�ݭO�i�̖>���ѓ��ޝ5�͚ͅ��ꐎ�]��A�ɓ��-�8�=;;�?������*(�/9`@�<]�Y>bٻ����=Z��� 	S�TU���!�:Kĩ�����9`�ڻ���@�oO�VK��v� ٹT�r��g���0��|�j�~v� ��a;��\���.y�,���6��?�`��:__	u�5c�D�G�}���Yt��T�$VC�r�'�F�l螬�[�nS�B)� :�!#%�+��e����� 1�.~��=-�6)z�Mk� 'X�Te=;@�a����	���˫k�x􆕫�{�n�~9����G}��<�6$,�f�	WZ[%��׹��\�^c�z�|�)��S�����x�Hm�����[$]z���Bl��p�R9��x_�sV�Ӥ��i|�]�щ�OZm�[����U�Zz�Ǐ�)�������n�*j�� ����m�R�����66�ݼ���S���Y�s1׳o�QF�s݇6����y{+����)D���s�/+P� �N������K��:^O�A}P���ꀏ�ޯ����޼�]���F��etg����GG�u_u�Qd^YY�zIC���g��� g����.l]�Fo����#����hWӸ��ǝ�;�$��?�S�\O�yVn8Ja2>PefͰ�\e)9�(˸��8�D���j�azz�
�E�-4�Jtn��Q��]��G�"g��$�?�@�s̺���?����/�xu���:8��S���|(ݥ"_�m�qR���	͸���
M��:,�v��3�QA�|���P�4�\4A�h�{�w�;�;j�]�47��.��X�e5�40NْS��U*����΄꥗q//a�XB�lx�X>�O%���|g�@��Y�\��=�{"fD��G�΀bM+�%���W�dS�ʕ�8z-��9Փm
��.mkm�~<��0�1]z�Fd��_��~s�*�#���B'����~��\::���I(W�+X@R
�jWjOAA_�RE�'5�w�*q����Țz���]�%����1M����7��[��s�[>����k�{:2ǄsH;J���"JmO�(W�'O����TSR�HsDڕ6'Q�Hך�Y�5�l.j��$����<:򮾈Nm_������O��T����0�0B:�$��[�E0���r�$�mz�pIIiR&����M���iڙ�~��W?����/ƆC���S����H��%-�)%+�
��K��U�is��ϊZ�X��q۹��&ݬCCC��w��ĳ��?wa��W�{��Z'�1����y��THGW#]��vM$�����6�Ji����
e���T��a(X���E�(�n:0��{P�����+"��g�6���@W�IU8ûg�1ѷ9:e�cf΢+�K�'�6�%"]��띢Lq������Z�H�EHx�؂�u��՛$;}թ���\A�S[>Y�[X��6����' K�t����W����Pz�P�.��T@��������+�,�R����ޑ�\�=׉=3Y�M�w%V�~�gs��Sj��O�Н��W�������X
z}�DA�V��"Q��g9�� �OǦ��s�ͣ��#>�֒���í�'b����{�}/����E�`bo>:|B���ρ�/�k�կ-.oV���SQ�ÿK�K���P�n)�It�P���ĺo<}�)IW�V;$h5m�����z)3��>�۩���C��8��s+XI�5cB�W�*U��/l������ze����k[��Eih�;n�vj���ߕ;Gm�$���-���u>���������s�~��y����p����� �8T"��!���7��?[���}��/�`��g;�9��-���Ō�|��k[;}C���O6�,\��iYJc���x-��j��������龧��U���
u��z.�8���'��p����%˜��`�{��K��-Z�y��ȇ�UznMY^G�&�yl���E�R��X�4���w�·��Α�`�A��8��fjE
t�.�}n��xFz4�������L�NE+��$�W��IC������\�j4>	�e��y�ݬԽ|�`-��1�s�d<������v1A��k��~����xJc�uYɃ�Ur"���%.8��@���90�g�D6]�*"8*Qhl#�����Xln���m�Xf�֩n�k��&���{N���ͫ3+��k&f��>B�&&E+�Sʓ�$�0�$&��(���ǯ����L
SfR�*���H��ERP3+���K�0ԇ^C�� �1'��K�#�MMM�3s���D�&=�i����?�^ЗyB���	�-*2��^]u��}���_��6c)�x���
_oŊ�T����&��X�����Sv�;|�?��W?��ϙ���_���_\��W׽�	IY�MbFb�����{�hZ��Ueܶe=��:G�C�z�d	[�Vcs�,Y;��l9?$
*�?��o�ϗ�����S�[�u�`+׹�\P�ӑ�N���b6�er_a;��#�ݺ�r��5����~��G�D��UV��6�~}��b�
n^e_%멃��4�^��z����Q���E�9� ˮ׆�Q�Ha�Q�K���:g�d���du�/e�׃\�/���[�M�C�V����;����ʾ�eԚmj��%�?Q)J��h�#��O����EM/�(%�J<��[e�ᢰ�֞�׾�*Ŕ�����d��-��?�P�f�i�6j���?�L��ea�fev{}�=������n�3R���y�[���n��kf{O���}3��;3">*D=ݶha<���_��>��9�
�l+((HZ�g�Z��j��>�m�%h�p�6Q��c}y�l׺�5AF�o,�B���#_�yv~�~H���?����vw�:F}�J�@��I��9�^���〇���$����r�٥�s�Qc�%��I����!;'~W0��UDe���ͽĆ��ӓ�QV��
�d#<�'�y3MJ�^�R���t��������}9J94�~�t��#��.��C$�3������g��nf��R�R�G��u�r��9f�F(Ok~.?�!�[oůlp~�������x|C�����Y��.�����=�uO�	������P������'�&�⻬m̈�sQJ�t���ݹ�I;}v?���?��?"�#���H�)zg���ݾpH��jS�1K ��V�P��=Hw�l6�O]1J��He��Z=2���tj���{κ�ǟ��7�v+ܔ-�BW[?��+'I���X��'�׼��>��9f��:�m�Aw|�x2�d.�`V��ĥA�យ�(�@_�%���.��,"�'�o�s�I�;0�[���1�y>�6oQ�U%���.���[�C�t�C�=�[dm��E)��-��#�*{�֖|(�L救�xUS����$�_�P8���[�;���iѩ˧'�Ӷ*ػPiB���'�-�|;�C���-�2��t�`prk��1��@�I�>�C�a~����k}�)om����v����Ob�P��דs�`\MIXw9w��6���#�K����&==�[s@w�,�U�9n0$�V\Μs�ۓ�{�b@1�[��?R�c����*u�OJ꘿��6+�El��۬�=@*W���҈����O����DY��y�Ċ��ʷ�����x�Ͱ{s����F*b�n]�����PtVn�+�9�����Ğ��S��rW���}~E�_�$+Vl{X�\w㪼�����xM��0"Xtu�b'�����z�uM��z��#V�>B��&�:)���ZZ��/<����D,�Dqf�ZJƅ���)��6C*�x�gVz�����Yԛ[������}�oH���=�A�G[/��8u�/�ۓ��ƶ�+������ ��]�|g�*y/�_K'`:�WfV����׉�a��P㇎����e�o����Q�S�R��(�

{����t��-iZny<R|�����Eov&�I�������.M<��6�n"
(i��?���9�����"G�}�[=e�8�Bt1ia�ma8�ͅ��\�F�_�v�z���ˇ�_:n#�O��S��s���Bh�[R��?m��:��o�?NH9!��Meke�ez�2�+6ce&��bg�3⳽��+�Ҍ��R�k�$/���~97��J�����߸�Е�s��L�������MGRz���~���vP�v����������)2A$�ӑ�n�ª����N5����r�����o{׸2�AŻ�I���tmy�O{�<�m-nxm*�#�,%�VUs�u1�_����>��U�V,:��=��ȱ��q,���_2<�"�V��#���#m.d3�:��Y^馻,tt�S�itt��=JV)�r�u��(=5�r>���C#L-����&߭�?�m��KܹKmh'�6,�sN�H����ҝ�m����{\T�Ua���������Gz)��u�D�
�?zq��Um#���N�kV>�g�Pm{%������%ir���b���f���C�|��J���׹�+U�m�v�6�Y�K���N�n%R�+�K��JS���Q����R�Dr,8�'ń�0��e��D�bj�*+	�&��2�������&x/�jdk����ֻU1��7ݼf6�[!�m���z]����C�����_#?��F���Iz�P�ܩ�j��C8vc���-o�EX�EU2}\6cd#"�w�%|�N�ן�������w�W��bB���޽?�;� �N�h��UYZ��������EM� ���թ�����_���AOؔQ���gO�~�wArT���MV,ݫ�W���,��(����<v�O�ɑ/K�w��)����I��E�t'��d4�"u��Q�1(�[hq��/6�ƴ��|���cbC�犍��8{_M�eդnz�L�A�a��� oL�K�.���Zn!��d3�_�(�0������_p�i0��;iӚ�!R�l�6j�༉�uH����ߗ�.���e9���u�%Ň[rž|S���%��~1Օ��{s���kf��sk��P�0aD���2_���/O�}�cYW7�z���J�(���e��K�ߑW���c7>n8��>��;}�|�G�]���;��.�[��O�������?��
�E'I�$9v)G�.��f�k�<u� �[Ju���q������Ys�VT�[H�Sf�to��i�P��/�9'Y��K��Ysi2�r���ٔ�]=rcX�.�9�)�\�L3BL��?��;���}���bAQ�bDE�"$4E�w�
� %��F���HPZ��!�"EP�z�PB�3W ��;��s�8����1₵�|��>�\s��|{f1��xx�3�|��x���3|O�iG�B�8�m���r�'�H�PG�ʱ۞�.I��Q��W�?�[+�&�Rb�`��+%�rK�x��}�_��.)ﯖ�A�9tj�̂肏�F㵂��y����1�4���O�,�J/.b�H�btuS\�\r�aolұ�q�艜�������`0U�T]R����R��N`�!���	�g�	i��jfƹHV_�6:�]~��z�3�2�g��GI nqR�#�Qg�2��C�2c�b���u
�eA
'��U4���eϸ-'|����E��+������?��/�k�?�D*c��[����ѥ���c�u=�Y���R���C�t� ��4���7$Q��J]Ӏ�6��)&a?]�d��`e�%/��.g�5fae�Dc,G+��~!A�2	-I�����r��������hJCʺYp����C��o�S��U�I�A�J C�E�^��/¨p�˅�.��u`��**P ?"z�/-2s!�y_���qE���ɶ��aݜoB��:bhQO֍�ṷ�A)�S��"����,�E4��;5�;Yr{�������dN$r��<� �%���K�i���N6d��w�}��x;�޹v�J)�Oo��q���h���~e4�P3��� 1�;PhL���F�j7�$Иk�loT�h(&�Ԥ���}O�g�ꨪ+��} ؑ���I��Q&��Oe犥���bG�mV���w4R���]꩞H��p,~;���q9����O]3^����R6���i@��<r�y��,�RW�
����:������G�{�vkn@�}8���*d�G��%t�[M4���0���xO{��<�IYf���#RE��u)�O�2��Q��o4�尿�%6�#�֭���>HJ�����
I/m����s�ט�s�1ӑ�|"D�U�˺
��(n�TF�7]��`���N�z�7i(���Sq�ֵs���X��҃���׿���{�K��K//,g�:j�1y` h��/��r4K�r�PM���m4~Fc�GISQF�㸨kB:�}�;�/@)ʛ��&fd��0����e�
�**ǷL��{+���x��8�h,,sA�=Sc;i�����#�&����J�W����#��U��0���n�y��V���N��w`x��6&��p#�i��z��<����*oi�o���_�w�_4A=������>"�^{��/vG���/���b_!����M`����+a�]��_Oz_��y��"�]�Sxy��G�������'"�Ul~3:!��+0rCc��R�N�7�r�/�T�r�&���T�괛�~��0����C�J�h�oZ�l��w�,��/���2χ�p�ع]��E��^��jcS��jR[ӄ�9�lK 6��.GT�l����v�1�N���R�g��չ̸��	 �_t�U�����,�7��Td�{�zg�#y�0���S��7�_���o�8�
���� �h�W����<弴�Y�R4kP�h����@f	D��=IIzq�ɋ#�_�P����6��2��
���W]����_��7�t�C�7�u��+�h����;�N�dN��?����@���F䩈Aޱ/���������|�f�ς��l��3B��~�ȋ!(�v�<[�D�n���AvW�/{��V�W����@C�<��y:C�3Q�2
�Q�"�So���=Gt�ܗ��2B���Z.��� T}����B����&�<��V��";��?c�4� �bW�]Ruv��Ի)��������ޓZ���IR�h"��g��^��?P���Q�ʗ�O����o�� 1���"R�_d����q�S�i�uɢ�{������N~�}�"�Z�X��W��u�Cc����{��-C��9�2ۍ�OǈK�e��}��\ 
�l�'/*ۊ�ك��w���&(G��[H�u�t���Ŧy�{�L�by��,���b��x�\�jSE*u�Rn��
��xI1������}"쾖@�U"r����A�=R0D�X��M/�$R���ݳ+ٓ 8�d[��d[j�}����#��T��^`ey�1(&!����9��2�H>Ewz��X�-M�tK����Oɇ����d��LN_p�Zv���v�nn!��ñ���^	��J �@a��Δj/�Z�V��j��8�~.]?���:�V$���)�Y3�l�a@Nk��$�r�z�a |Dws��zv��r�cs�g�
��oQ��J!3���K��+g���Q�]���oZ�[{�� ����{���M�s��|��\'~�݄v��'�Jy(����Uc��e���i����_db��B!�;sW�{�v���x����5�aU��2�}�&������Pz˩��� ����۾*oh�]{p�co��z?
�;��IC=�	��	������ {����Z7
�Fr��뤘'Lh	����fC .c�DQB�Tcm�'����'N[�LD%&���
SĔo{��k��>�9=�0u��JWJ�eI��=��z}@����Hr��Ձ
5��8��c����4�c�/,J5�A	wk�����Gd��9���� 
�Ի/�%�@q����2t��=�󏦅����f�8��Hl�&��n��.OWX���s]UV��^���9�z�z��~�F%����IK�}�d��	�P	es��/��L��d�We)\5�z�v�ґ��´�c�A��� k���<���~�W�����Ꙏ�f4�9�1]�$}��c���p�ƲT��I��|B�k�YM}�༃"r��ɀҁ�a}�""wc�7H�p�KzQV���9z?��(��joi�΍�sW�f�%,�N����j��O�I��O��������)M?D'��y�c'�ͩ�s*\ Ƹ���>�'?�t���2��H�G�$c� ()p~�N��V��`nc�R'�3��D��$��k�P��^���&&�EJ%��CH5�%�V��ӡ�E��c1Ά�٠���2=���%ÅrdJ�����3���)t\��C�Q���8 ���a�,� X~��^�@v=�
�����f���I{�}��D���o�L�\��P�#f}����9-�EG�c>����� 9ʋD�E׹�nD��3�c׻�
P��j�~�X_��sP�*��!��YU&25aL��r�eD"���~�U���鹯S3�p<���P-w� ���~�������(��Oɇ�k��U��:��C�~%�L�0������2�������N]��<�i-�9��;ya��94%]�.2 ���D���P��r�Ʊ�etN�S��q�Zɮ?�Ez6�����9�
����6��b�'2�_��������+kH���|�5!k��hV�xƧ(Ue����S9��MO�Q2wUYbV�T�2�k[�[���R�90�Ѡ0��P�~-�v�&c?�ߐ:U1<�-�8��*��$W2*ZΌ��9�
��.�k�������w��Y��M& #D�¥,��q_�^e���2c�s?\��4�?`��\$x+h��Ty��/��6�I�"��Y�5w��D]�8И���}���l��Z����}+���Uf9v%�����2ФQ��̔�0��t�:TT�,���h)[������=�y��c�� v�����QM{~�h�KLKoG�P����*ui��T��lU����ʎ'z�]�0��0J��B����Ť����ZǤ(DJy���a���)��RoM�o�w��(gP�U�6W�5bC�ث�XȰY�m��</�ܷ�:�O�z�NS���ې�Y�g�B�QPR-lK�Bi��Z'��z�=�r�3V6���V]���\Ա�C�y��!�fI���kH��>j��o�u�#�4az-	���p)�\�ei����V�5��O'����eȞ�Ъ�������.��	��������d=Lο�x��2��i��/�����	*.�������IJ�\�K	�bD��N(��N_֡��U��!+%=�f�k �m炱����B�0hԠ��Y#,{�]��4�0\ )wx�������^�Ѓ�fZrHx�*S�e�kŞ䰃,�Z�P�s1!mǷ��g�Hر��1�����PL�޺LN��R+A�R�a�� ����s��`��g�����z2���"�-�afy�bh��,�o�h�YZ��b.��]��{����x�1��k��0�3;@�n��FOf到� ��v���W�86jy�I-;�3����~����g8��������8k����+��_9��_�=���Y��|�H5��=;�n�SX�����dGt����i5�@8�Ж�ިX���g}�캈��h�R|����E��J/� y=V���aĮܵ���x�=���y:4?�T��O�����kǎ�[x��Ž1���pw_:�q6	�迓���#��]��ݗf��&��IE����^���B�aMK0D�#K���2�1�k0�ٔ�A_U4sb�U��*6��M%BW����Y�4N�.�	���m�_�b+��q_Ķ\pq|�N�Ǿ菮��z�T�.�	������ݴ&�UO��k�=�_�AEu꿪x��%�P�,s���$�p�y�E��V�0�oe�b�oPm	��v��?Έ��V����^e���:�������%��5���8sC\@�L�\�t·\v�1�|j���>ij)�`>W+���`�k�D��-S\%����M��eC�)���c�x��%���Fn���R,'���a��-�`v�#�3}��3Z\�Gk�e1�a�l����gT����>���q��n�x�

	1��{�3�{�]��9{K��	�@��
���M��O�/L���M���ύl�.E�bS�� �H���9jQKDJ�ne�U_NX�}��2����cc�����r�r1b	X^^.~2��>T���=��ʵ�\����L�ݯo�-T�DˊM��ފ�^i��&���\�Da�'A�$K2u���mֶJ��-12&&��1�7���/e`��?�>�S�e�Q�Y�U�V��%8�_z�1�����U�|T���ux7,���������j�F�WB����E�����OK�������?��?��������g�حm����g2+��8���#(�+1-�H��8>B�B�UB��2�hהPB��3����19�E�;����}E�7>yO�R;w/]�'���K��h���>�\}�v����/ND���(�r�4��R��r�N$C���T �m,|��v���R4L���фM�:�>~�����7ω�4�q��n(.�֣[���պz}���Ob��w�-g٤�c�����Xf��q��J�i������=�!�����tg�;�����A��c�l��y`�]e�R/:`\k"YT�|hX�/B̈́4�����jω���Z���m���&�ض�����[Ô��ݯ���z����ve*�'�w�^,����N,�~�{���AW~���� ������OĖܓ;Q��ЉC�.3�/�+�lj��1�ؖ2<����A%�/����Z�~A|e8�D��LWqZ-�y+���Q��/�1����Au�:_9�3�!9{�b�d����婱�@�lG��n�
��7;r;���Z�IԾGl,3�H��?�!���O�C��Y��Í�oO0hL5m��~T혐�|�5�nT��q�[�����YY��l����O��}�6���t@��O�Z���P o�����g����gr��i��ӟ�n�?���D_/ ���D���zg�Z�idzD�/�u&�/�:?��Ոsē�����hr�,q���y�c���αo�ln����fb�����;�����XqJ�L��?��`4�_�@%�_��������m?�%�
*^
lGh��[�T/��}�_-t-|��x��2ڸ(��Mb���r�����OxiA��s��M�:�G	��ߓ�
:���mL�IO�{�I�?H��tR��
�6Z�G�s�	�Lm2#aY`s^��C�6�i�Gy;����U|��γ��Y$K�����6�j�=��Or~�/�����S���%s�hFOX����c���x� U�����?��g��I1�4g,;�K��#��05�՜)�To�"B{Y��Gzs3j�ú�?��[�6�u�]�Y�9����Ũ�a?���me�]]��94�9܅F-�B_��h\_����G東/_'�i�[�x�)�rn�Mͻ�r�X�2�4�q��%�/�f�y�jH�"�Mz�
J���l������lR��_�=6�茺5i&g�LB*uCg��0�&D�hY�S��l}��VA@��D����>�ͥ@���T~s�}��މ�tx���p���q�!�R�٩7Ʉ��J�7���n�Ն��S�~��8��aR������m֬�b�~&E�����rq�g�C���}u�W�j&j�O�;��D������zr��o��H�(�|������il�;�-��}��w�D�i�X��,���W��mwB�ܜ1�9e��[�^�h��蟏$�k&
g��YD��X�"��q���18�z�@,��▓4�E���܉K��uV�T���N;-f��f��oC��IO��[>�+�a�t����U��iA�D�[E[��jh��ƣ�ԋ,/w�寐BZ����GJ�5z[��>�TR�r�i�U�>6�1E��ǳ��(���כd�:�)'a�J�V��s��jN!	��:{!h`k�x�$
��"U�m�ơh.[V��X����ΚM
:f v�����rS��6���w�-ھ�/[�/jJ.1�GJw6L�R�RUWf�T���6�����X��u��<�����T�9����XB�2�Gٙ��؅Q�U��
$� ��7����@ qY�l��/o%�D�P����X~�Dw��h��w}"(�q�\ջ+n��-HǋhLfxv $?��Й���D����1��Fev���.L̀��A�,�!�����=>,b��AO�Z:c��}�M�^��1+�U�ՙ[�RE��g��ތ�~vS��[��T���7J��l��.���fqȷ�2-*�iRC�{�i�1�������8��<��Д+_�v�E'!�A,���e���ȎL`�J�\���5f�¯����/t1�?�R_+��+"�2�7�s`�ki��}u�.��.��K�b>+e|���&}[�h����V@�א�p՜�	����.x��z����i��&_��\�n =��.Q¯�1�OCe6�}6]l�A����ͨ<�d��1�p���bS��u��	;�kS����������������W�1���mX#'�`�r,����Q!Ĉ	{�W��Ȱ��.�)�$ljz�˗��y��S��l���1{(a|╰f��w����ܛ�3�p���~l(�rK��)��N�l�mձ�K������R�h�3�`��a�����U�rub��0�!�O�+%��}�̊.ݠ��B��[�(�F��(Lz/�n��T��2'���Phk��$ ˽����!�n�ܯ5"Ν�fLpXq$º͙�ax��v��ծ�~�|�V�9òc��'?(��
ԭ̱�*�8N���6l)�=9�B�0>=9�3H�V�R?�z�%�K5s$7΃�I�B�fj���V�N=���L,raAӼ�
�x�a#S��
����q�Hi��Չ���߀p�Kq��#?��vm��LX]���=ej��bi�l�N8l�ϕ}�q|8&|[�?H�Ŧ�G�N=#�A�Y,�OK�u�x��ᤸa*���?�"�mH<�m�s$�)��9�ߑE7�����B�Y��S>��?ĝn�-��A|�O��r�>!�dN�L��?�^�<�t�#m�G~(\�+�E�x<�~.�<{Ǳ)��K��O :?T"}D���p�\��y�q�T�o���ʛ�ג����shu�W�'U�s������5K��<h�}[sL¸T���hB�Z(���N�D��Q���T�N
hξs��s���/��;�&��^�}�Z�a���3̨�o��=�L�
�{ç�*���۱Ŗ<�u�����%�MTM�Z=�g�4�!W�P�)S"z��H�{^ϓg���1,ŚI��'ɩeia���nB�v�-_�<��T;* �}�#�M���͒ח�}�?�Iռn& ��>����4P.4��h��@I�![w��9���^�`��_CD�uޖ�~��70� ��!&�2���k��}!�~�I>C��᛫��gyv�D��I�q����m���[y�ՒϮ.f��5ka9�,%��t���x��(0��C�*+",��=����0CW� "Ӫ��ݮ�����Ge�Y���q|��g�A=\v6݋���N��<cm�RۺN�ٳ��)C�pͺAݞ ���[�V���S��N�!�~����e��_�a����>���z`�WW�+
d�C��!���~����%��� f�VG�(�Wˤ$�/
O�2.f���V��W��}�k�Eԏ���UgD:n@��a��~:���6h�ϯk�GuZ╎��t5�T,Tcy��������Q���m����=k��4��9q�*3�_H��q��c;��٦��,m����(�
�|,s���e�
����2��X8�0H��Ɉ�KHƦd ��jvSVU�G~���CZ��eXE���@U�{ٔԫdP��<��~}
��k�V�釟����d�3�|{��{
��?��x��ti�o�l9��3{����̏���R��vp�,�Cy��#�\��{���6�e&ˇN}�ed�춭t��.��u�6�K�N�4 ^�*fTw���U��u�詚��)�*���<�s�����F5Mҵ�܈ j�-;�h��~	�OR۔T�)'������Q�khL����"#7M�u���Hi�ڹ'c��=+:?��z����U��Po����.)��ʵ3�<�<j;=%�Z���+�P8hFup˼<o*1��$�q�*plUPFZf4M���j�,q ��26�b�+�@�a��[~ئ�c�m�U�R_?tt������c��!LB��9h�D��je.�!����%���-����M�����{��t\��V3�j�S#{�'�v�5G�<�> ��u�%=K'N@�o��^�_��&�9�>҅R���x���B�js�04���O��@qҫ��Ɠ���J����7��Ep����	��HY�\�j��Wq�^��_�����|�ٜEZGvu�^�yڻ=���4���Z��[Ъ�w������D�� e᱊�=%N~)���zji,(�~�N�t.4�G��M4����|�\8�$�VR*�f$9LX���:�4�0���Dn���R~���B{_��̰�� 8Pc������:fͣtU��NUULps��(�|��w�`��[|�!%���~��aA�p
���΋nE��[l t�cU��׹�;��ih+�y�@�����N��[~qPϥeY≰��
�8�Yc�$&�؜�9�kj�2�K�O�SP?���T��C��'P;�sD�1G�n�QiIr+�cU.�B.,'���uU����nb�\\Z*r�� �Oi���
h��0[���Pă���WI)����F�4`�n���L��Oƿ}�t#!ͧц��}l!����Ufc����^m_��Q�����@���� D[�N����#A4M�-RO�Y��7`yO��D��(���6�-�F���HbR��|b����
��+��g �,K��:8p}����7?��0��]˩MGa&cu��Ft(�j�䇞������qL�ӝ�t�ya���d��V�`lh����Vg/=�́��$(���= ���2X�k�o�)P6��ޠ�7i�-�+>�ϧ��a��o�.�����Y�i�����R�U�Olŵ�N@�kG���0Az�^(����XE���?��zS~+v*�j()&e�(�A�����nn!�>��j*)0#�s������a7�x� ������̉����[��eC�I�xq�T-SIY�崩c������;fR����sm>۔H_zo��_`u@_D������Ƣyކ6�QfH��޸��TS��|#띺ܹjt[~�o�Y�R
�Nu
a�Tj�� ����K.q�w�&��粼(��p�N��O'� ��Le�'˾ڔ���eϦe[��������#ݓ��Y�t�UieP�t~�'_�B�B�S������	x}z��)�U�8i�Nd(h΀
1������sQ3U/��"ʽ�L^�d�7�K��(����˄���&#�� 7��m�g=ס6��^*����`>��
��V�9�̷���&/ٿ�![��[��w�!:	���t��ƚi5I\4�E�9����d�n���$�'�ʗ:Y�bퟺ1�l��5�y��ħl���˻4�JW!UNZm�mu�?�� �(�JV�Rp8�#'\
��,�6��Hf�SF���x��]Cg�����R��*hIjK�Z�̰N�W�@�I�z̷�H�b�⍟�V	+Q�-�e/��U��g�������;�H'��e^ӱa� �i uK�_�~�B�H�y4��{�y��� ?�q./�u�_[e#�R�#`:�E�|�a+�~^�R�@4���� �D�=:�WPc�Ҕ���ضP�y�TA��n�h�S���a�qu�t˝�*m7��N�\:䷥d���+J�C�Pa�*\I:tM��.9�y��r��ko��	iG�^�7�w�N"�ԏ����}f��j�Y,4Pz�3`��A/��m�
����ގ�� ubL摫OK�q�dq�J�CT�/$玲����Mb�g���
͡�YR��/���/mTd`7�n��d��xP�)Q�W���ؐ�wo�����9ض�\ ���wS�:Xji%ᤲ�X��-C��wÌ�:�e��U(߁����%�?��#�y�iׅB�� G�Β��|�`��T�TGR2�{��j�-���`�h����:��ȧ�.���C������P�˗�׍���}�~��xt|l�Y�9���c�!L�cIs�Ҳ0�;�[��2���4��������gQ�����s��1G���D��>MR��۱9LS��`����f�|���	�Lʓ�UG;��;@�q^�4����w�|��+I�.�Ѧ`'�ZͰ�g���$@,PXn#�-��蠖H��	b�:�[H�}��^���pQ6��������G9�w�*�`{3yh��^+�8)����l�.����/�a)\�]�*�1���'��h�i�A�SM�X� �vt�@�%�k)fa�Fux�kt"1?1�u��pV��Η'���Ql{�Vڷ6^�&�B�[����g����+�F��}w'���	e��*�~ЌY�5������z�Wf1�uy�E��s���?��6���XB:���  �uA+���7�����+G�T��a�J�+69��y���!*�ѽ���I�J�Of�a(�\"�͡�&q��F�p��>}�jf�H���|�18U��DfbOl���1�(A�H�����V69�G�����k9���?�mh3����~�� �R�zM��	� x�k ����@����GuѺO�D2t��m�8k�t��mщT�Ԏ,�p����5ӎ�<�mX�ba��6tT`��J$r�v7M�(��m����"�:�����u�a�2��{�tSt�|"6����EM���9�-s�3��lE�+����P�],��=��@�%��e0Q:�~gށVtr�i_�IKmQ�̪�C���OȌ6"o������X�uF�zeB\N��G�D#�c�V�|�S�C��m�'��P�'���7��u�C�2T]�)�~yX�R��ab�x#A�Y�؄�����Ne���Z�.����8��?М~�m�8�?���:�їc\�r���\V
�إ��	�5�^���m\v÷#4�_	�Eԍ5	�Z`i9�G�Q�I����t�o��d\�i�
k�C�����b��M�iuI7@���8?�*g)�<u�����6�p��G���<=�� 4xg�ywM5��%7��4ԋ�1�(���)tnO%8�d���d�l`<�d�4��!�;"-e^bh�:W�s��۔3�h�e.�L���������!��LN�*u_r�oR#����z�9  �(��r����<���Dv"��)k���~ꑺ6����PE;�Qr����q��L!�ۏ���Ay���H��A_�)��&�l��w����I�M'���PQ��f��\�XN@o[��<�
��.����"JіD����bX��:�`}�n�+����.wծ����"I��m�0��®pZ`�u'�8ծ�i%1�+�[�'�@-C�Z�����e<�T8�1E����X�����]��u�4�P"�!M��k�����{�n�]f�	��ֱn��ׯ�Y��"�*�>���6Ƈ��D >x:�tbLї&����A�8>���gh��vf$�j�����itYQ�ϙC꼶�F?�zkZu�r��Nӳak��k��,����d����v�h�"���{u��bϽ��������Q���!�����Yi�)����~�l(�ӛP�[�"��[lr�Cy/�F�+ؤ��6�sJ���;vN�Ilz�ne����U����[�	�[V��)��#�ޛ�ei}NQ���B���\"m}zNw���`�Ƥˢ��ո����>{w�/�� �,�J��]����C6vLUp�p��A�z��ą����^[T]F���ͣ�S�M7J+��T
+3������p���u�t[	���|agjG�|Lh��{С��xoa]��"�J�Do������;9�<۽]󳶞�Kȡ;;���.��z�ۄm������UO�DR���[_p��\��Z��љ�3c�*S>�XyjtU�É�Z!��|sɃЯ��<�1#����L%�Q���Ȧ�iR<�@n��uwJ���V��t7�dt}�v'�(u���3���;ەߘ���LUn1宧�����26����W��Q��"�s2���x�׈�	qƽ���e\������7������l���;}T���,L�_���ᰲՊv�<���u��u���JHZ���S�Q������."�]�FK}Ɯ���P�C�%��35�V��#�(Ƕ�ve��ں����%j�T��o�������\�C���$Of���=�2Bݠ���PO#)�z8i���D������X��Z�&$c�������V�����6�,옍�0��U
8�57ֳ��?��N�� +�-��	��4��R��l����`�/(�mU��6/"	d~�ݾ%��rw�왱6@ҫ���L-���B�͔�jM�F��ׄ�˼�ݎ�'��]{IR�5�xam�Ys�4���͢j���3H2� S�6���p��[n�J�B���sl{`�6�9r�J�-11��EҚ/\\q�1�u���C?{��pS
�xr��7_-����dn.	Ҙ���U�8/�:�l'��d��U�Fw�er��J���?��يl��P&}b	��YX%i���fz�,�������.������Y3�sU�%�>�j7��Hh5W~'6�)��Kuh
�N&�����{/M������C�2�"����PE#��=i(����b�d��W�Z��/kG���
�9+9�a���H/�����*Z@d�즐�v╽�PDy��/�a��5s���m7(&)�!SAz��wy/_����{g�=�	\X��e5�xA~�Qw�S�����O��p��`�����B#oV�V��R-����(3�읜��EE�{+�z��Ā|��k]WT.��ӧ��k,ct@b~���g�WPA���m��/ވ�����Z�T����mb�h�lx��3�:��*v���6"�s&
�bǆ�C��Y����f��}��F(�v��v���{����,�������|�SKcoίz_o"G>I���5��хNc�Cw��0	�bAm՟_�����$h�[Fr��{�MB�i�oVlͷ#,p��w#�h,���<c���H���x��M�}���]~�z~�e��>�@��;�>&3�k�u��T*f�bt�^�#�xv��b����bE~z<�O�©e��"���Y[oM�F~��˸�j2VY��N�bMx��l�Wmkh�Dm���p���� ��!��{a4僥}� g��Pg��j��)^�b32�a��w�t��M�03q',HLL	H�\[b:�h(��zR\���;}LS1�b�Cp�U��\Ut�bݤ�B��EU��:͖�kQ������5�e
����?`���S����8(�<BV����C���ǝ�z�d�5���&_��	�t|4�łH���f�Ά&^��k���U"~� Շ���X�ʅc��i���Z���i��Z�R�\�f�g�]�>��O�~0hEsg�ě\ߦ��S��Z����A�]fD��h��������o�����d|ǔT1���H�7p���b^����_���$��SS�$;��,���v��ɤ��G/s�=;��t���,�<zVP>=�J��Z~������1{�yܻ�4�VyGւ�|"�J��lqo�� ���.��Ü'�Տ�ֹ����]�h�i�������4{�Dp8�Z�<]b���.{y��1j�����F(��T4O�d�3u���s���%w/��L��ֳ����[u�\x�����m��*���C�pYp4��gB��](�B�?�t��C�y5%6���0��чt���a����db�QgT<F-�쮍58ii[�&����o��H?;ĪE$����TX�73����l��ɴ�W�V쁪�����O�|����:�6j#�V����4�Q��9�{�j%S��Vl܉=�(��j_|�x�VO�P�G�feK�_MGy�q\��3o�.���"����Q[��j+q�W���ZU�S�	�^��M�"ի��{�T�c�3��������	sKn��%�BP����+{.�	��4�ύD�L�<���CΕ`x��^����Jr�};��reIƄwO@��{6�v�R�G���-��>���*6#��u�c�=��c {�̈Ǎ=���}u��Խ�z�����tͭy���t�׌�ߒ{�T����,��kW�����T���C�aIIg�Z��s�$[X�b��tv*+�qB"M<ͯ����V,�OTfK~ݻޟ��z��N�ŊE�CJpe��(�̱�/HL�O������O'�[/.��҆���+h���nqOav�#a��rۍo�zgg�MMz<Ή������e�(w���4���UT$�Z9�nʾ�C�Gk��:*vRC�/��n�?aR=���>s�����1pS������ݕ��<�g������;	�rm��%,���K*	���J��mX*�w�Rǂ^�q�����R޸�{�<EH�H�����7�[s;Kh�tW�?q�O��C��'G�W���Sy�t�k�z>lq�A����Yk����,�]�)�\�1��D���z4�%N�$���m�m�$�A���x<8��m�Ɍ�ʔ	14�i�3���?��pp+w��碌@��X��t��\�{$��Q���wf���obΥJ�=Z�z�)�!�d���ѶB3C9��g�#ḡog��cd_S>��'��w���n��dvv� C�m��%=@���R5X%�ٕ����=9�E�ШV(��=�� ����+g�Sc�b��+��.���-a�x{y��.��ɟ�:��Qm�'r�#5=+�V��l�H�(���@�ѮԨ%��m�b���ߥf��W	䳦W64
eu,��Us�7/rsSc�WGƍ�����,8_4.�p��G�%҆��~��9��6>��,R %`���]N�V�F��HA`��Q�8��~s���ߝk۵�Ru��A��k���q1N����5ImX$hv\��uD��ԑV�_�2a�ۺ�I�Iw�32���L���x3��H6��������2ȣ[c���~ye���`Hp7󺣜q- =Ȓ9>s�zH�t6~&E˹.�%��Ҩ/c�U�E5V^D�a��u���N�K�7�Y������3�w9þ��ߔ�u���C���2w�c���]�fK�J��Dk�oV���n�i��v����g�I�춳��H[����<����2h��>����*_��r!��˜=�}��k���?�Lx>?r1w�A=�*f�]�i��+���?��Z�j-=�[��6[K�s�ۿ�'*$�{��J4���T�Hx�i��写��v;xs�G��3P�9l����+��C!���^G+�y��Q��!�2yZj0�M{��$�==Á� ��߁�T�&���|��kC����'��S����Tڸ��"^zjB��@��i�u u�$En5U���� "Pu2-o=��������g�j��M��*[�6���l`�Qj� �Cc��^��/�昑(�v��S�d2Q�U�wa���ϿjP�i�`��HÇ֍j��Q�G��fY�zZ�R�(-3��8�xX���tQ��B��k�{�U%�iq�7z��Bh��g
���o������k= �u�Qc��S��4�� �c�0AN�5W�� Yz5�g�T5h$���h4bq�d���1Z��%z��i.c�:�uC&���Dzz$�E�`�߾g���4�?�l��w�]�o�@���/fkeU�{�yL��['G�5`ԅBCӞ3�8a��,W��9�$0�W^	|3���E�7���8ػmX�����[��ڰ��'��e@@ ������3�,gf�dV[k�HQq���y��� �[g�A�l�XU����6�:��_�Pb�3��k�g��[���D��p��o�NlPU<ن��](;g̾a�g`<Ei,q��?c�� Y�م�V�@^e
Xy��Z* WZT�4�[�!~����O S({�po2�}��bD0��J��CO��Ae�laV�"�so�JBl��U"�%��b�-+�6%�/��j�\d�ӳ���t��3�����_����D��� �Yx�0˝��]	�R���m��R���᠒-��������w���V��yk��-o���Ox���ڊ��a��QU�E�'��oC(��v����RjB�v�?���#��x'�Wa�\mљ���e ,W1X�Y.彏�Y��I�f��XE��͞�tW��RgU]
*���|o����w��N��j�g�-�H�:���'���=�_W�MX�i��sת�ً1VQ\c).��K���[��rwm��_\�k�[D����$~}�������H}�3+�K't>�O��a=l������.=UyA�	Ya��tSt�R��Y�;W���[4�&ZՠǛ��)�	���cr�@ݻ?ݑ���ͯiX����$���=Y
���^�q�]c�����>7v�����y�Q�J7�E������?S�-�^���B���]�M,m+��F�+A��[�].N����ȯwIow|(�Di��@Ttt��ґ����:�+��=P�L$�H'�!����莧h��A^�۩�yս���/횑S�w�Q�R��bc Nʘ�3���P�j�rϒ"��X��R���?�s�h
Ι�Ӯ���[}�;)����5@���6�m��2�$����r�������z��Ǳ@���.E�Ai�IEB	)I�R�F:d��iF:��r�{�{��������7�f-����>{��y�9 �-�Ij�_����a� Z�f�4͉����[#�7��P;���;��:s,R���X���l V������~O��߷�����x.�l�&��9�����=;���JBݟ�7�V]�MD�Ql�ت�Ab`�̭-�7M�R��E�e�?.��v������`��\%��$iq�&h�|0��a��u�g�ڨ��9��T4���aK��`�����cqNx{U��[�ۚ>����?���&[1zQ�����h��A��I�V����D<b��_ ���e�� �1:�_���Z/&�)�u��2�!��������{��b���,&99��'��쭿{V:Ŭd���G��z�g�P�8������b��	�8Ku����q�Q�fc�ȉVq`�7�Ȫ^�>�4a�IV��l9��ut�B��Q��v(_��q���ܼAn^`'N�S��4��4��-����ku9�Ȳ�����S�p&1��*V�����J�V�Pkh�㟡��n��hۼ*e
��#_��UW��a*����3�0�еd��"�c�q�?"��Ā�6��x�:�3���'�q��A����X�ٕ��y�Zt[�hQX`7�[��nC\S�2��ە���N?��+Z!ۊ;$$@(�w�}�`R�X�Qj�;��=(�=:v��(�Q#FGk�a(�sjx��֢������HL65�I�-j5��N���̠�%J,����ϛ6r���ѡ�%^H�6�Mq�޼���1��6���H{Nɖ@U`��"���NL&|��2{�Y����G=�c�!^�S�F�<��(*�[re🡶���,��Q�����p}u�ͳ��N
�w�~|�ڋn�j���,�j�Np�*�S��o�KY��fS���u�T6�#w��wvܷ�I��ȑ�i(��Z�<�0�'��7l^M����]]�'�z2�O9h���\��0�k#d�R������fqUR�,j����ΆoT>���I�D�ƒAm4f��$�V9)��f�j�=��A�vo�Ǘ���O���5�Z��<�\¤�&z���/F��V��h��9��	�Ye��Q7,h�VreG��  2Z⇇�
q�_�
n����#��gf���'�P���hB@㝂�Ҟ��ő�X��Mݡ*�7v{�l����dY����WQ/����ɓ	V�����"�r����w]�O���;�J���v�L].������կ�2c���X
L�ťƄ���5���u謪��@��|0��B����?�T���7��
8��#����^`}�شN�8�a��'�����B���'#E�/vuJ~���+޼���hމ�IIv������e	U๕����a�ǍU�A�#L�&j���,:�<]#Z�HB��>_���y"/����m?M�I݉s�W�d�&Z�	EA�1��^�w�[d�w/m:�o'��Jl�G��o ��T�0ub2U�ٌ�6���B�P���Pm��T��H>�����i�`�SB7�"f1��M��,b�U�+�_�\G*Z'K:Sse=�0�S��l��˸V��5:���r���C%�+������hV�iND݆Dw�K��t�C=TU�E�(�!}�8�k��@[M�=��"��"���Z��T�dr���_9̿�C)ƫ	�5�9�����x�����ɻ�gs�%��!`�IN��9 <0x�~����s�oŏuD�Bύ��:����������.%��G��K���E���=]�0�b��FU\M����dj�7�qo�I�46l��z{vVr�m�jBC��؞Í�;��h�y��̔Dv�4��L��x�wc�V����d�0dX��z� �&��s	0��{~w� +]���Ҷ��������Sd���Yԯ�����E�>o­	-���K c�}� xd �V��'L������ŷj5X�������q�yk�TV���7����=K��X�L����p�U�D��P��g�~>��8��M�q���q��?GM�$5'�?��7�?'Qd�s���Γ<!��9����9��q�������~��E�9*"�y4��y^�9��X�o�>F.֭�nӛW�p#~m=�Ճ�5ޭ�m$��ͦ|�fX*�����P
b���Q�E>��)׈7VJ|�O֟5r �R�DY-���ah�6$�V��\�9�^��0X��,!/�� [� �I�nl�t���b	@f�����*m�s
JPP�xOO�xl��@fQ�G �̻Uo9�GrN5"_��P]!�G�,�;xhKU�z0kE���*/�-��]� �Sw�^��������q�����S?���+:	�[Q[���%mL����'ۛ��W7���lp����b�_!��i��H�U_�/�1\pX91�� ��̻�����o�'�ȴ�%[Ͳ�jy\<w*9��i��릦��P��?x����()�����A�A8[��}ۨ�P�=���xf'����.���>f� �0�,�Q&�����3��`�'02z.'�b["	�q7g��&o}�sV�Z�J�JW�Qb�*:��A/�����[K���:��n���vf�sദ��q���m�&yfQ�'��/{"��_ϻQ��#�d�'�.�ʘ;��)I�|�q�8���jG��A�2C�6�xz�Ǭn�/6���Tq��l��~Y,
���`p���s<|Y��4��/��p��Q\_�9�ԠJ��~�:Ҙ"�ԗZW�����\��Rn�M?�j\f�N��@��5�i�w���hw�C\���!���rM����,9��b�>c�S���O	h���m�7tWY�΅��T���0pH��	��b�s�mA���շ�|$K���A}����R.��uK�ʀc0�J����*��
i��t4Eq�� `�4�*����kc�X��T9MM���2��w|�����6���ۨ�4��l�(E|��|�Q�p��w��ab��ˆ[o��*9iͶEg�[u��>3!�'a���T���D}� �����āo�5ޫe��:f3�\H	��?QD�ɸ���Ccկ{��<M������� ��T�n0nBh�"��~	�~gc��Т����}]��NS�C9q�����[����Bڂ�������ӛ����	dS�Nv�c�ĉ�3ZƑ����<�tt�B���f�X��=������������Nb�Y�Flt�J=0�+w��#@�h}ON���I��i�A�.N����x�|�*sT�`�i]M]*�@ᚻaú:�Ƌ赡���ޢ��b���e`��> U1yN1�	QL��}��?���<8@��J.7 ُ�r�hH�P�����H�\�͈́Q��o�xbF/ب�����>��g�=��o�mfM#Y\�n��>� �!�ie��K7�5F�߄�cJ1�K1+����9����xZ���.I$uJO-]�b�ȮȠ��ǘc�!v�3uV��4nJ������'�[Op=Z�Ԋ���(��waD��{����/�W��MN^��jQ]����}5_`���Qf��\�1�}�̼Zc�ևM��s�M5��|��ߢ�B��4�1�{L�4eE:�TT�(r�h^�KQ�0���0���F�m����l�����|z.�m�Kʞl�_��]�_��r�T�.{��H�kq��u���07�b6%�(@(��C��%��kO�R#J�}�;�67��a|���1;���)�#��&�l��6�߽�\1+�$&'{�Q�T?/c��`.�� ��"aM�2�,E��ĸ@4/��(���0��UYcn)/�f�������,�'�&��~~�{ɫ�ǹ����Z���FO�*�����􌾭��[�zs�N[�4u/<��wG$�ߗ81�9`���gh�j�Z"��i*��� �M�ʁg"��\MF�9!�N�HG	 �d�m����Q穡�'�]b������4� ��|����髟���Ft��$��
>��S'��[+�JI$�a�v�����U2���k�����nn~�KU+���I� H���h(y_`vO�� P�ؕ��V�.؄R�5<(1B��@������0��t� f�?�?�݊�r��@?����ZIh\
�$T�h�ߛ��)Q UX���)�E������T�1(���͍#U]�)t������`@$�z32��1k8�c��Gzq�Kߣ�0��b��#���ƹZ�>o9w]ii�F��8$ܞ���<�)q����5)']�y�u=A\7~�t�6[#�,�Q��v���u('A�s+)~�&j�Z@����=̇ޅ�'vtts6�шNC��Z�b�9��zu�G6��|W�f�z�hN��^ڐ�O��e�F�s97�gH%��:�?���Ǌ�i�V�TW�`��"Z�:��c�r�A�v4��,߁~�i�<�-g����lo�x���0��-:ij,��3n���#�/�G1���DPK�� K+������p0���>��a���f���^���/K��yR�
�z�2PLJ7k���2�\�MY�ԧ�1�G50��U�{����4Z���V�M/�;��&V��J��M��gݤ�S�l�t�s�xeL�C�Y>m礴;:�����fͥ3����� d��9}��w�7��坼�b]ыm����y����.V��V�&oϗru&���]��"r�w��=�gR������;���}ȃϬ�~w}��7 [$niOK-�Sբ��4ɻ1zG��]�b��7x�Ž�y��L�����G�����01S4kg���Y��/��q�N���?� 8dx+��^��-�{<���n�����oeaF�6��ۍ�7�����-Ƈ��}|?��\����n�ږ�h�YJ��x��B|$�~�ҵ�uMT��8Bީ�<���57�^yQX!jI5��pIx�j77����_�0�&��FM�XS팧,uC�:;��Lm#=��ބ"fS����s *�@aˠ���w����u_'h1�=q	sDA���� m�k}�_�pÝE�t�#��j601�F&�(I�~. ��g�9���e���z9�8�ٷ@�h'��S�	W�2�ă/e���D�%i^�����o��%K1�����?�b�� ���� Zuy�~�Ƽ>zv�=�'؎��;O������K�u�������]�p̐��z,�ѓ>�	7`Wn��b�ЧML��*���\��'���A/-N��}�	mx��V�6�)�K��ŃEr�&��l&�K���J������~��3fE󘕔x�^zT�E�-�AO�ߓ~FC?^�\R�H�����|UOr���~T�3�h��6�+�jxѽ�U�����@��8�B��6�,��3�Ɵ��v��H��xn'�JB�O�'�Ę��9%�p�����m�����#j����a��I��Q�@�
�t�[�Q��J�B�V`�Tc:i�H�k����Ȋ�Ut�]�6w��fP�6(L%x��"[��.�nxOꙡ��x�L)#z_��J@z�"��o3����y�N|=4����6#�-Y1h���-Ɖ�����S����y�$U��N8Յwd�w�����Wt!��d��7X������85���TrȦ�SC�OFurw�\/���º��j��䐊e@I]w^b�L`�J5:,b{KE�w�5��Ou���=�Ŀ�hױ[��q~)N[H���$��&mD{����'L�ml��>#�-ٝ��T�-s��&�imhV��/q���y6U���P&If�-W��y����1+�c�"��v��͇'o[<�Q�D��j X�n.�ޫ���;j���R�y\�������bo͡i<�㙙�5D�IfUý������_{��g&�8�OܺǱ����8�֣0*�m�1 �<��M6Hn{��mm�h�S�ng���3�M�臚%�MSP�y,��JV���a�kEl�E��R�s�NZ�	,��U�Tr���:e'lЉ��9Q��%
6�r����AuT_>Z��y�SmX+�k�H�#�ٗ'�t�PB��kr���9����MGG����w�f�~�����������g�'��8��x؍'l2�S�ѭ�1N�9q��輮��6���<����N��R�鈴�貨�[$��1<q���If_2�d ��z��l�I_���r�
bw��;|8�^�����m^{�
�MI|譮���tmM==+��� ���J�n]��F�Zy�ƥy@:1Mr����v)���<�ml�D��љM��^��5����B�[}�\#��,��������S�^5L6=�)�
'�ɜ'm*&\1|��ik4&�ְ;s
Us�{�������sM.TN4�?p3���>ps��vm�F�����ܓ���ֻ�X����h�(z���r�q��r?�-h:���u����e�r�h�'{�x��W�b�5bD?x�yvݕ���7����6���r��r�C�w�
} �<
�}��M�3���r{�����~�i���T��D��5�5Y��(�·ר���Ȉ���H��8�V��Ό����"T��Dc�1���2�M\B~�:��Wkir2@���zz� �^Ao���m��D�;�qX2�� ���1U[cw#��;χ��:8C�9Fl[�7t��	�N@��Z� �ߒ��y<c-�l��%��5cR�#�L���'�`��9-���8�	��

A�D�X?�9���o��z"�H��v�Y��;�r1T)����x�s������ϻ¯�c�����3�qF'����֦ㄪ	x����Hp����n�]KTo{�`��h�|Tdj�}"��|6@9;H|����r2���9�F�����5������w�����1�~� 8���~�!�Δ��h��9۽�+rz�������~���Kѽ�G���s,�e�Q@,gݝc˵̯�u0yQ �j)ʺ�mZ��3����Mg�o9����+1����O��C�����H��i쬌�,����Ha�.6i���M����W���Q
��) /']1uC�^�v:�狜����R�6L�/}5��V�걠K̩�`Ô�	�C�|�����fy�6!?��zjV���oe&���އQߋ�G�g�1�@Ϩ��[S�Lʡ�ۑf��p��V��@�b�)�RQ�fY/gn�I�[�^�c]�o��Ɉ@9�"߳^���SQT`�@��͏'-Z\�����Na�&�iV�d�t:�<�X�O���:����z�܎�c�7#e��(��D�Z�7]�^E!�(U%�k�]�����^�2k���L��݂J�~���d�N�&e4߼��e���	d��&z*�,�.;��;���K	�v��T��H� A�_���Y��m~�S����%ߢ\�w1=׫���9[P�0����_F�;�;�¯���V�fsY8hޕK_W�N��iy8����iEl���m#�	cgg`A����"���(߲��[>��~P���$����5Z��x�rDn�:�$�O#pz\�͞�=^�'v"P �,��W�?��Ǵ�o����Ы�xٕd�w���vn�?K��nc,K~�U��9˸���Ǵy��(�
2�W���:a���ɉD���^��k�?�r��Z��A����>�fi�������f�װ%���@.3���հ�[�)����:�>7LX��!�Wy�h����Ф�����WG�܋�� �g��l���|ܿل�I��|��������%���|�e�9��җ[N&�܂�	馻C�<@S�(^�y5�+2Pe/3ԟ�3�"��B��Sˤ&KȞX�cz\_����N>���p�Q��ɞ\sӮd6��6���-�/S
�4�2A~�v�_����*L��{�pT)%r���c �Է_�x(d�����a�لQ����Ozuub�9w���L����,iz=U	��Ͷ��x�B��08
���Ezs�s�����q=|�/�T�� O@��`t�"�y1����x��iqJ��Go�pz#�|��y8F~�JE�X�j��|�S��x{	���M����R�Q�<�f��9p���NS��J:FڻKKo����궏�D<g�{�ތZh�i�����ܐMZ�[�b�bmI����6��q����!7��k��n�߹��Pr����3-NvswX<�V�������V_�~�g�U�r����-��/W��S�`�M%y��}YnL���-��J��Ř93g�����"��89��B�I|�]\���Ʃ:�C|��D=VǍ�T���D�������7�2�j�$���ظ�$�:m��?z��#�.���~�B�gyު�Hh���=`{>��;�w�}��p..�����������i�������G�Q'٢�t�W�Х��>����Ŝ��ϋM�����'cD�'�SI�W&�]��p�f/��������iEw�a�?|��!�i4̞xkg%�2[p�aC�9f!�i��m��`*}��BQȂ�ݸ����
��~�B�e�YCD%�o����={V��E�2C�QuW�y��s�$������ٛX���G��^K=sȟw��⬝�Vf�Qo}Tc�x���ˏޕ��[�ߥ��%�?��~F&�>O��9I��U�HYVo1�Y�z�_|:���'T饕U߱���ϱ�&��|�v!�(/�G鏦IG��ŉ���u��m���zu\�~�{Ѡ��Q���ǯڍ}HBY	�����Q,�N�#6�G��L����C�<�����k�Rͣ� �ȭ��	9��1�r�i�G� ���-63�5�BBiB��ת�5G��^�"	�c�ܸ�~��C�k��.�^��U4�c�A���f���� v�d�(cw�ۢ��v�V��᠑���4O I����r4���2%&��%|*�?�MqΊ|���y8�G�]_`��K�K꿎��w�@�vN���]�Y��R�����hoa���YV?�T=�K�>/$�/Ù��ɔ��v@	�j�Ps�㙙�W_w~��B5!`o�U�����ʆ[�W��l��'>�3�K�D>N������sD��oUi�L,�����a���Kۿf�p�P(�dW�|S���AV4��ŀ�pV���Z��fO����H��E���J�v?m��^0�M6"�"T��*��6��%�$ �H�?�$���h[��,c�(�i8O%)^���͸�gXE��8�v@UGy-�~�V�y���&7�4�-U�����r$c�=�����?n�\)ɗ�<y�G5�ZI��c��[��0g���n�����r�z�H����(I�5��+F6�����fL�{�6��ȥ3;�&���S|9u�n2�Yy[]�y)I��1�F�O�7�o��O�t�&q���_���T��� �m�5֭�t�f��u��ȳ�?J��b��%9����CՋ�#���F��d�O 7z��~��3l&H�%��L,��̈�{^ȿ��s}KZ����һ㏃�c�e�-��&!}�W�'	�[�}I�u�>ú2i�=S��Y��:,my�=-�V�c�d�&��%�BT^����.���<1~@>�0��7�V�S�[`���vQ���.x0��g"B����#�)��
������T?-�*�?w�ut��L�Q�6ʕ'OԾ��|myjg;�vv^!U�h���nr��x��_���է�V�
�����N�o�d�G�e���O���9IdW�+}�rsT���M��q�
�yY^�Y��n�ˏ�ik�_|�-������JZ�z��×x�{���R�E���\%؉7���0�҄%c
�&�Mby��3];��O���XX��_�k�3��C�_�o��Ng��K�/q��d���yDr�r�P�w�MR�{�+���w�y/ݹ}r�O��js}��[�����eޠ+�vB(���Gx&|V^8�dX�T�P'�E�����M�0�Z�
�U¼uN���� �&w���M�$-�{K�z�[��iiߘ��Sr.����{�p�]؅�[ͽ��%1ߊ�ӱ!|��r:3�T������d{c�1�-yY���6��EQ�L�S�(O��h�]e��P	T��׶��ӛ��*�ʾ.+��#�t���`U�����F��[̯�Y`��5$�����~�E�{�ho~ >9�Rs�P� ��X
k�m�����DSv!��~I&�
	?���eܥ��Q���;���ƥk���VĪ;L���!q�������E�gV"Y�>�>\؝�+A7�m��c�(r���N���
7��!���%\.�<(�R����r �A,�*��C<�ϣf2䈙�,gf���r�[�IJ:HnT)Ʌ{��E�D �Ő��27>"X�j�6yYN�y!�@W��Ȗ����#ܕ$�(}�6O��e^�rԞ�z��^�D�c4�:L�t��� \�l]5n5�>E�o�iB�p7^��&��&�u�êby��ѓt�� �ͣW��# �����ȷmM�+jI�Q�(C�>+�lgf���u�f��(*KsR�_^yA}j��;��}}k��u����$jB'r̔�g��|[A�J�9�6�?�؍��*b�.���1���$��$<����2�i�ՒS�d���rN\�Nugi��'[���wށk�S��tzu{ �m���/�k��>�d�\��^��!=�൵�`��'���d��Z]Y�_�Ժ�[o��}5�S��#�)����H��`��8`c*4b��|����1�}{��].��Z���#��퐪��)1��z�?Vױf�K�|D`�K9�V:6��Df��o���}�b��6��5S�ȅ�~�s�Wb�$���q�¨�BSS�����W\����X�;��[��wX�Ωuo���8�a�¬G�;�A����d�v]2��9Ju�)�~�A?�b��S�6+�RqH�5���
��Q�>�
|6Z�Å��
�z���	òq�>"�w��0�p����:O�Q�R�/�ll�nG1\q�c{6�U�&��1���V�%{�q�L��y�5*��&�G��y�,��Z�M���C¾,C����~#�`m�[�C��߃c�[�V��i|k�m���y:�j��v7�i����gI^Je�(	n&,)X6����<�o��Fy�;�$�NNO��΍r>rt5ͩ%�V�T�|��=�4��d���C�{�O�����0�]��O���Aa���8�_���H�Kl������ֆC�_��R"�R\��p@���3=���N���I$S�s'�.����2�/ ����L_�>�1
(6�w�;TH؝�=6}��<'�Ē��rT mj˾F�:��[a�)k�3j_XVM2{ؔ���-{^Ha�LL{�fΖ�Ő ��U##���ѝcr�O�p)��g#�<�=�"d�������{�?�ǹ$^ύ�l��~E�G�����mm�����?#킛�AFePH8r�f�f�-wG��[xM1�̅�x����<!�d�;��%����v�H��麪�	.����C�bD�L�ԧ֋k��b���5g�2;{w�A�
ۚ9yy�&&&'�kk��i���}��P'߼�w馟�O�z}Np}��i {�����AZS����|�SW%�h��x�˗��<����{6:���nsb�5�JvT��Ųq+[a���$�L<��'
�V��W_	mI�oZ���d�\���^�9p�����#��?�I����u�2T�Q}*�!aU���y��������G���/�w�F���a�U���[��_<��6���u�m^>������ޜ�|)�>��Ҥ��Ȍ���_�g1<]K�)�A�����}�Bdy2�GYYY�a�Q
x���������ce��gB���K�����=b	�).��5�z���(�2V3-���s��\���P����ڿuv�k�h��M����q�-)���8��!��a�O� ���ͪ58 m�� ɶ�u=p�4��vnu���~�G|�"�<�?�T@�'!��݈��5SE�S�2�&��K�����Oe��H��/Ï���캹�z�/Z"�4�_����L2NEE�������G~��{o����k�-4ב�a�-,���j�T/�0X�D+�W��O6�=x��[Yt-�
JH�2/5!��٘i��sޖ�aV�`b��O�����K!��d hn��ş�
��%�%�V8D���;��F|N���p����Uc��_�Fy��9	v]5@������m�w���#�N�u�*I?�SܷY�$+H��Þ7(>te:d@�;��x��A��M⼐�T�'�j�r�0�E�.#i�΂���O��)��F��xٞ#�~�N�H�_m�${R%h����^��=���g j�a�a�4�؅��bHc��{�ۧ�f��ك&��� �χFF�ǌi�nc��"��Ӂo&+_�����Ud�G�Pg�c�dg^X��9d0�Z�=Kkg�;�߻|A��Ҩp����'G��@���w��RU�lWU �Aȳ�S���`�;,�X��[7�m4��'���w7=�/
�7iP��5�R1��-O�V����w"Ք��S�nM�?S�K=�?�!-T�*�#�\�S=�wf���^F�9]���|T���k!|Oy�f�����[�暽p�N���[:�\��%3��i�8��$�-)^Jp1)�N��C�����y�=�b� ��6HY(C�z辶�5��}Ն���p��7��0V뎹GN���xn�D��3�^H�٦�m���f��z���.Ei6�}���'"�
AYO��W�p��Ԫ+���������v��K7Kn��*���_�£ׯ�'�L�5��gv���Y�$����P��P���Y}���w�z>�7	�Zm�Ql�n��D������@��m��yQ1$)r�	��iS�m���9� do�f�5��/V����chȊ��w�Ą8��}.����@�������6����-�4�)�eh8�� ����}�'.q|��]em�Y�T��k�5�'-�ؕ=Hf�ȕ�3j�R��_�/g�딾�J6��#I�}�@��d����p�y�K�wq}������j�g1��k����A$b��$��0D��ȈVye�|O�e, ��6ާT(�7�L���������2$2�����W�? �8*n�
}�u�@�%���'��b�����H�j��G<�
�J�������o�D���r��1�z	��x��,�(+ߐ��;�`{����t���a�s����g1�c�+7��;w��WH����ݮ�A���A��𮡜�h�[0��		x>�5�f��v�K�D���~�g���d kw�o�
�Y��wܬ���m�}Z�)���+-�X۴i�>��G�z�/'5$��E�v{>m�[r��j8�*6ۓ�M>z),pteZSgw�z��˵�%O�{� p�R���į4ֶn��d�'�v��������I��dݛBYP���-9t+�K��~X>dV �6� �1������Eڐ��Q�/�/��hia���EuFs�6�ttt\/(��@�5�/~�E�sA�d%�B�^j`pp���6�P�����Az�래a�> l�V��	�um���/�k�>u/_�UK��YL�	���H�m�5^�Q��7��q����K�S�$�ϝ-H��M������N�ǙE�k�7"�u����ȕ뎓����J�
\�9�x�E0s�5���UQV�m���ꕳ�Gm�#(
�-I��A��o��eݬT��a<z��1����%o���p��sh�w ���6t�{FF��G����$��i����w�ES[�5�{�b�:��;E
��V�����-�J��G���y�`�I^,i*� �� 2���3T\��Dy����OX>���eH���A����[J�`="`:s��)��q+��r��,���Q�W���i|P8�0՝;�#l����-.�N�u\���'��ld	4����եߋ�s+h��x�ro"b�}�e���@������Z�Nc"oJ���A�7��_�����0���[���1���_L!/��Y�MGH�	��䛳� ��Q"��vdo�{�h����$u�Q�@.|_x%��W�q�{w�qN�I~�hM�1����O���d2�r����C����A��M���Jb[41~:F�T���R�i$�Td�����=(�`)��{�
��G����\�]T�:@�����r��^����aPY�LͲ�c�އ�����<�}<<t*xQC����#�!���r<:\Rc��;W,*����X?X�x���<�Pc%.�r�]�F�;^�.�Ǒx��b=}77]�U�y���
n������'�Ӱ�wx�R'؟؋�h���vc�f��Q<����	!fn4`c5̑�$��ʳ��id�$Wɖz��^m]�p(w�GX�\\@�1��b��k�7��MuB�hZ��_qcأ����e��>Qm�DiL�������f��L���=UL �N|�4RgV�������`�8���Ʈ�K+��/y_��7޷{�A՚�����e�:'Eg�ϑ)��"��S��>�tYt`x�"0j�!?-�����V����@�HǄ��x�s�S�ٽH�����4�#2��m��:��j$�J��L��L�oݽ�����"�v��� O+�Դ��My�ɦ���|\�v���q��b�x"��FtW���nA<�7�4��^��]�N�ߨ�(�Ҵ�I��������wn�̧6i�i�pu�.��M�V��I`P�08��H��>�(2+|>��=���;��7��n���N��8[��,�:��ੲ�M����2�6W�g�X�j� ܬ�C���Z�b�s�ъ!��g{ko�����";$r�?�f ~��\�6�u*�JSSS�ƞqbr�İŧ �j�<=BT��U�thb��N���ņN�#�����GL
?ˋ����t�W=/�:n���Ȫ B(7����7���a_�W��&�06�c�p,Ҫ�Za���v��oF}���
�Lqw���)�:2�QZ��9:6�_[[{�`L�~1�,�K?�tw��&AymdB�cfd��R�S���pݦgN�?�x7��P�~�Ɓ+d?�ɥf�|ڂU�}1����SY����5���턦�������W��f�F�jFx����!����tL�G��W�*�PavB�Ѿ�{�U�g��d�(���Svf��n*����뽫ч���F�-O�ǆ! KtKt�n��/M�/�~կ\��#�<����y9��n�f�~��M_�P�η��~oL\ϸ�߫?ݪ�f��v������%��	�d#��I�ɛ��1!MV6�>�Iyԙ�8n蔼�VdV��
$^5��G��������n:!jp������+�r���'��I|����RK�O)�2��>[�4ҼE/���)W�/���}���2�L��
¢
x����]O��8�Pm��Ɏ�\�J��P�8R��S��bp��Kx�^�=^S���6���?j2[�D��Y�eˑ����Q%��_�����g�'��y@)1������6
��xT�x��ݱ~�D/�	��KjW�Rzܻ$��J���j���(�yg$c�n;��Bf��'��1���s�ͦe-��T���8׽�S��������H�gc���5��I_S	a�K<���e(���T�"�{�=?8?�k��G�Ee��,�rI
f�lm��Q�d�;��~���+F���ƪ�Z5|]�N+.��2\A��e|K;�K� w�r.���C��<�a?~SHI�W�Sp}$�J/����p.u�,C�fW*Z;i�(�{���p��ȳ�-K�&��� .��)[>==�FH�u�h%"c��$����y����-yړ�-�@[�k���=�oiy��sf������y�-�z�=:~��:㱧\,JN��;�/�WQQ�sz��CЦ���`��3����{����#Ň>L�{�f<y���_q�����3�x)O��[<I@�D}�z_�4��w����;���[H}�U�.�ۼP�}5e��wjX��&�1#+,DG���ڄK�d��2�ζx�1L��%]����������q����z~�a�R�1;���}��ϩh�Df?}n�����Q':�v��R��)"��p.�q1i�	ͩ��b�J���&N���D	�M![�����~���L�t���a\pZ�h������{���D���!x"�+Ap�(�pY�<�e���<y�dd����9�	�l7���=4U�e@h����#��w��DSs���df^qژE;��YY}��r���u_IL���a�g}q�E���#R%������}8�F�g��|�W����4�ЁbU^̜azf��X��苷Dw���OE�ʏPG�����#�'�v���O�����e�v�2w�����G�ҫ�t����Y�Tf�:MY(uq�<jr�tG��$΂�}��he���f�\��v.�+eK��Ǎ��Tu�G�Q�Oyq�fIC�(�L��x�o,���)��x RA�ٷ���RU��$�^�Hr� pD,���}�%�[�(0w�+p��,f��3^pӪm��E��^M����J]���ݏ�w�Z�ͫo���)C�ٵ
0u�����]�4���~>��A><<<Vb��p�Ly˄��|�t8 ��ՑlG�Rin0������)%�uB-(���ב���#���t��Ru�|���+L�1;��h�ӪaCRg����뫴^����wno2�P�V���MI��k���8�q�"�N��u��sb��bp�}4������yv�}L�$�[��'��O5o.��z��R���65RhYӒѮ|���~2"�o�\h�_>P�_���i[���2�p�\��@��b "�MJ�� ��jU��s��P	�(Y�ʏ�M�)��)���]{1����ڹ��J.M;�7o�c_�X�`_'����Pޛ�&�u񥮎*==ݟ��R�hz}�m@Q0EUWW����/P3�s�p\^��Y[�Y��A��Q
2&H��� (T-�)+9ާ�TB�����SQ��j��~33�G�������1�,����;l��ᛓ�ׇB�~�Ҩ�͗�+�WP��y/��v����Y#�5�.���Ol��Ll�ҡ;B�,2G��܆C�%�0��f���6������S�	/�;CY89Sm���>+�T���'q]R'r�R�$�o�}��[",�s��� }�����U��;���w^�E,p��HuHF�ܲ��+ϸ赁�F�ߢ����<pJ���m�83)��l�9C�]��Y�L�@[I`R�w�uk'��pe��z�E�ϭ��Qb�~+[z_9�癭�?������>���"!�"H��J���-!�ҍHwKH�t��đ.��Н����{���ُ�zԳb�9�kͽ��ח�!����V����&��}�v8T��Rr[/ϴ��f �������]>k�mAro�@Y��IO�f|�L��x�c����s��\��č����Ɲޙ������
��L�oW�{'���2an��ܝ^��XQ����@��ի�I�0=�$hu|qe��
GFN����>��Ņ;;;[�T�=>s�H���7w���P93yId�AB.��9&�_G(�3P�!!X�dX_�*��|s8T���W�N6$<��L��������4�@��N�=NW~�𹽿�Ә��X{#���'�����͟d%��~��	[���R)2/�P֎�Uib��ob
9z�Aٹ���\k���;9���8���׍Π�����n�`���&=���O!��v.�U^ẫm�!v�w�Ls�q��,l����FM�1�w ���@Q2yab5�oo�iݔMRI�r�}�3��'�f%�U�'&N���u- C���3���<�XJ�ڵr��;1����굧�Ѕ�>t}�������퇯#K��P��@�F��Kh�dߥ0���fs��Oɥ#�5*�f%�L�Ϙ&�|�����y��_�F�#��݀������e._H4�Qt���
~~�N�v���?��#��%�w���g�%$)u��3%.Җ���@�>�2�@��ǀdIBBB)e�{��~��e�-�-%-�ee�J�&�%5ޒQ�&R�>0�����ru��_\^�Dw8���h́��>��\�z��U�"�oL�ޘ(����s��&"m�F�v�/LZa/輏"L��ƆzB���11�
�O�ϥޢ�ƚ8y��H�|u�r8d�Z{F�������ؼg���'�S�[�J���m�ɷi:�<z����wJ�@̱���$�v�����u0g�wg�(���d�Eȋ�(CF|�<��Ȝ#pK�.�?�[������(뭟��Ò�b;��I��8�4��YC`� �F��� y�椻or<�LyĶ������X�H<A9�B,	�b��of��߽ٮ����{�E�d�[���վ�����s�׷{�>� E�Nm5ʞ�b����X�`��U=2��J��o�gd_~��}T�k�B�y	�H��R��Q/jy�Szv�G�_�P��"l��cض���/�{#@�e�E
� �{�>M��[��v�`<# 䖺����[l�@s����he}����P�f�7QCwߟr=8މ�{�p�S���;����+�Y�o���F8"������F}w��3��(�I����H��S���MR�-�,Y�P�h<}�ڮ3����8��}>�s��xG���Pkzz쌡Ȉ�����|�t���������n�CE_D|�ˠ��0�HE�u����$�>z2RJ4��bX���jd[����ǝ{�=wC'�����JlP���AZ}W�����E�i�ǔ�B��ժ��� 5�J�6i̓�b�,w�W��.k�><�U�pj���7�B<R�ጿ) DMMMw�����Hd@ɗ�`[�P�[|bo���g��F�?� ��`�������FZPwD�}��m�pm��WzǄ����DPP�߻w-�����1���>�
���Ύ�q�5x��֣��D����"ы�i������p'��s�a��#��,~�P���f������)�%H�5)���ޮ�ܨ˜\UE�H��>j�޺��>>M7���rX/j�d��e��7�x=.�V߆��J�7O�A"�޶����tqqQj'�4�� <�2)����Ν;l���,�&��x��tyKC��0������]�?\�8̌��r>F4�Ӭ-�H�Y>Ackkk���5x$�j`]�X�M{b0|""Q��`@)����00R�����ݿu�Z�/T�b�aaZ��W�y������Y�=W�[0�v�lSz�_�ZL�].F���1j��0H'��::���T�����d��������Z%/�?�\���e�৑�U��U���9���B�f9��}K��?Q���c>��z�����p����7��@�Q*۸��(��������B����A-=}}�@s�@�P]=��X��oy���9S:�1�ߢ�ˀ�l1���Xd����x " �/}: 聓����B|G''�хg�dd��Id>c��]�����j�L����k��.�iK܄Y�Ӡ�ِQ)��o�����m!w��wD��rpPj��f��P$�3R߽	xRz��H1k4�ߠ.�h>!�'��P�e���:�]��M��5�;�o������.�A)�^	C�6�����<ߔ��W�iyG��=�=S4�3เ�n�ˑ��G�0���XqG�VF��R6,��G�.��X��0;����Բ���i���f��7`�u�M˜������[��)�g��xcĴ��`�A�o{j++	&��7�}i7y���(�q��$N�!�RPP�n��D]D �ϽD���"51����C�bbbr����f;�ԯ���*V��.�	�����X��������r25��;hfL���v1����i,����Y9��8�O���0Hw��_�� ''װ��8�������f���"`����t*%wy�z�6֪�g
[H�66,�yn�0��a�^�i�FA��|tt4�i/b��>��|��w
��jA��,��>����)����1!ǃ؋�����|�*(���}�ؼ~�ĕ�K�ϳM��^�Ǒ��0qOL�O�w'���&����w?� D�T���%9��-�F��G >����߃��0_�b���� �gb�c��.�7H�1`500x-.�����+k�xu��U����{����ρ5���'����Q
?�咈�J�NG�ﱿ@�~Y��@WqYb*=a"~sũ�Yy��w�:� ���&�8@������c�7c9�T �ѽ�{(*'��<�Rw�g!'����uy�(���ej��^l�������5gG+��$����^B	��s��)����\-��e,�������Q��uH�����@�c:��`aQ�!�|<���>���e�s��)�T��Jnl���h���񝬬����yZ�9 !�YY�>p����������@��@�zUK�p_^^�ַ4eUiф�j���/>L�����7��c~�yI͢���?0%� _�8j��z������`���;H�\���DX=b�X	;>���<���; �f~�&ce8?�Z|�Xcy�e������>y�Qq0�o9b������l�d����V��QdH21�`Ee + �h@�� ��IZw_8:u��<_R�4a��M��Ұ��m2R����uQgA�z�&�ņc- n����W��Џ��U��{r�e��S�c�!��X=�k�Oo����|ҶQ��/��*u����ycu��(j.����B�����AxC���1y	Ւ���M>����_G���i&0<�����C#���Nŗ3�=^e�Tj���tݍ���b���$2������x��
�<��
2-�*���lox��z�(5'5D�V(��V��֗��EG�W1����m��Дs&H�Y6��)]��G)��g�?�J�'������6v�!h$�̼</06�u��	v�H�\݆���"CM�|�Y}�.C͟*�k�2M�Z(4��4/0PO�W���
ƎQ?6��<`PdT��A�4�>U/�����:,���v��1��7s�=���~(&��활*,,��#��M��_.%T��R���Cו�"wk���p�~�@s
�l�H��� �W��m3eu�.���)!�F�N�ޱʑO�=Z�4�[R>�X�_��5��tDZ9��,����ga;�� ӗ�}�9;'N�K4?����OǇ& ��1BĞ�t��xzz������r�h�.T,$:113��u�~+	~a]�+�6\W�τ��?���.��~@ $���ڍ�Sd��J�,Y&r�Rڰn���ŵ`#�'%����������(5	�J�^�F�Je&k��cn��ǈry!ɫWB��ˆ^�%qv/�{��A�&d���Q0�8��= t��Nw��(�mm��)X�;FE�YyjY�K�/�)K ,%�I�>(ۇ�Q��de=��U�S8Y�?�U�S�:^�?������W-p����z���>c��Qxz0�.w��^�4vU&����H��	�����{=`&��ʣ""�KKq�ѕc�y4j���	�(1�Hf��vO7�~��َ9��*UZ�=�}p��`ra���������]�i�_1F��i �-m�I�</YY?766�"#9e���7,Y��<���P��38��(&�����P���M��M���6�k��s��}@������%�eC��αo��Y1g�������:�
:��
�n�F�j,Q������ E���$Q2��azs_J^��B)o0w��b��}W"�����Ì��*Ԏ����W�z��	
��h�#-�9.�>��م���l�q
m*c�+y` �a�<����V$| �`}��MF.3��`(�7`�n�bs����.Ƕ���� ��Om)���z��Y�K�&���4�O.��txr��eP�t�1@�6f�')!��(� p!��B�Pʷ��)|?FLq�^�������bl�a�U�6ݟzQ���xӉNk�St�/A�	?ොq�g�?�5������k���G���5 h�a(�izF>�>g���>8��?0P8&!�  !!a�ؘsC���_�D�����Ȱ\�R`���	����-���U�V�(j
��|c1��9��m��{a<85g�ݷ���OL�+_���N�[7 ى~eN��C1���н�?`p����G���p��M�H=�¦U͛��E��~��C���� �e������5K�X>�U��C:�G� / 5b�ajJk�U��2EEE}��b�͢�=��ꠊ�J P@ ���qC��!��Q����b���n��p(s��bN��멙l�WD�(=rt��Y�^��V�]��s��w=�/��� 芑�?����IW�h�_��	&��}���{�S`����Ot�⺇.�tѻ,�w^V��EY��<�;F�L ����#���;�;��֏C�t�sz.��YY-�8{Р5��nw���k�Aƥ*5۝���sQ7`����7��K�o�Q\A�2�
�~���{��-1B���F|Y���S;��~�C�_?J�yt�Hq
j�S<5س�&��_����{���Ǌ�O����ȅ�JJ�g>�����Jr�
��V�Y�S �AG�y�ݽ	�w�N��'T��f��cu��$��Ey�+/,� ����OK����(Pݕ�+o��d9�DTD���uS>����I{�Iz"��H�&�TҒY(���d8�*�\�"yjNz��-"\�sk�9��E8:�O��E�`�s|���ԅ	V�NY����,�m��?cK�`�QX�ڒUu-�Iܿ(w
`���}3�g6�^��}��U�	��h�^L{1�xף%�7^�yV~\�iD~���6$|�fT�����J���}�[�y�5�� ��O�f�-�%a�wv%T�Bf�_U�I�j���Ė���a�����
A���~XU7k7����ZW���� @W�#�x� ^�S�`	�z�>))�(Hk����ӧ�� ����L�핿/TB!���0��H�L4d6��	��i �V5��<�Zq@�%G3����xϰ�r��9x\f6��ȕ��W�ߣ4n-aU�r��+�}��q3ff�o��n���j7�����4f;j
&՝������o�O��UU~���A�E��c��˿�/+9�i��'�#����ӗ. ȗF��O�+)��_�V(���=��-/O��E�y����UT�Ć#Z�?���~`#� ����(x5�F3?�xBvp��@� 8�x�xV�� �#*@0!���d
Y�P���*�<�SU��4�̗�D�hR�U��W���v������g,��;�K�#Z�d��s�Y���^:r�{O���^�/Ŭ��9U�HX=y-�}�q�Ipt��m��u��rJ�K�xq©B�ʐ�/�:�r[��f,;���TtYvJ���	D���f�ܮ#���΢���-s��F��no�b��b�y�ʺ8y�����g5�b����jdb޵Ї-ɕ,��=��ő�4�e���Ԝc����/\�NM�׎�~�Xw���?N�Ǌ��e����@j�t�Ç9��"�A-i��Ɔ�D�#C��:��ĖٞHz��u�����ݜ��b$��F^?#|Ѩ��Ja%����)��#���uU*�YŹ�<� ��@Ǖ]Y^�	jyG��iϤ#�[��=�kB�gaGs�z�2������������ǯC����pͳ"����˓ob���k�p�� ���')�_��������\8c�Zh��p�;i�@.� �����V��`�&�k��1�8hw��ƥg���n�ӆ�1�n�;�y�϶:���� ̭J�c��_C��@pyκ�_k�U�(bp�t|r��F��f�6///5p��9�׭���X�뵷��I�ۉ����W�Wh|�b9n6?���p̪;E�����}�/{��UޢK�L&��&r/�I��B�tw1�r�Z�u��>��T�ecc�@�_��˪�R��c67/p�
K�,+��U��(�⡅�|� <=�<�u�I����S�_�M���D�"W5]^�
k��Q0���i4������>�劙my��9+�r���	�:N{=,�'�4m�$�{Z2�Y<&}���X�������cƋ��ݳ�n����0?�|<y^ɨ� ���mbbB�E<�G�X�+�=>��6:x/mAMʐ��i?y)?Y2�I=r�I.e�B���lIN��Ą 0�ʥ��/�^@�߾���-�pn����t
��;E�_W9��@4��71�IK'/�ep�?h���cq.JS�9������.*Þ�#�d���V\���6d.���si��ۆa�R����c���jf����-��"��#PPQID�ie�A�S�lU��W�D}�����i<���kg�/ق��(��/�*�=s��ڮ�������B�"s���z�M��/:��ggS���m	Z��=]�|5����J�Er��2���>�u�S���ٍ¹H�����7+�\Ը-�B����j����˖rr���a�,.vK����� ��=?���, �z)+#qF��-6�2� ��8��-��>W^e]�=��h�b��w]�,�w�-}�8V�q������v+*
���>I�<��X+��������d_X��L��6�hf
G9�����ŉH2>W�E�w�\�sC���
وI-�� b�+ ���"x*+��9jftMT�Va���4>���tc�g�kW�V>��
��ֲF���C�(d<�a:jd` ńOl)fk[���)����D�=�/^(���vq�ǃ�x�+���}A^���ҥ�ei
;E��"�|K*�)��˻^�����R�zjQ�baa����,���o�܅i�����]\N��41�}�&0���Zɯ&n�t�^8��Ө������u�!H��cV��5["�ey�����о��?>�}e����w��T�/��'�C��-�rG���O�Zf�ΎVl �c�<:^$�w�X%7�l���y�k`�R���]O��1RZ5�J.�(QaRTTF{�H̳�����څ���^�ac���ngʑ�A�P%zib���qP���ά�Ĥ�~�%��R�N��?0���=�>ZLeF��@$IaR\\ �2f����	�Ň��AC�M�P�5�k��ui�iFԵ�����.����٧1JfI�Ne��3�*��J��s���~��ھ��VDY������O�H����Y9`����u%_���UTLg�{>#*��"�o\^L�t:1)�`$ @
���:9qI�� ��1����H�Pk�aSJ|U276�[)��_]5��헥������e(���ة����x���E+]@W����VT��0��E�3 Q7 ����1(n�o��QVj��/G�=@�&���}�/l�����6�Om�T[�țZ�W,� |
D/��7�J�k6��X�_� Hs�{�YF�%�o�����W�f��)8����r�^�� a�T��4ŕ�
¡�6�G���
W�Uۀ�D"�x�9+�,��)|�nUc���?,���4X�eU��䝜�
4�8�k����|����#xv����%0b_��І��y�j"����4
�L���RVV�xv���ӷ�$7�i{���
�N؈w�4Љ^�E_F�����e���m�Ћ6Z��7�F
rs�=1y��Փ��!�`A�����r��hFr_���nU퓘���{^�Vwl�0֔���426&�@��)y�3퇚2��vL>\��d��bBbs:,*Pƽ��������V���7�ǖ�B���E3������R=ǥ��_�ж~����!��m�Z�Ҳ2#--�_g������ �:3
�
�N�Ow5�Kњ�YY}��GfUK�\�G'�q������݌5Q�%?Yj�NC�@���*�񔍌����"�e�,��T��2�8D�K���w�ხv��㸼�f���=@d������:f��G���d�%X�22qwNA�v^A�$dwCì��u4I�K���[o��hH�ք���§`�\(���t�A�ոu�(B�)���XN���4���`b���Cȏ���G��H8mŠ���S�ת���N%Sh�ԯ���~�ӣ�޼��ap�I=�&sA�"���ĵ�CG�,��u�z2��)<�PV�]��IWU0�n�tS=�1���&m�.�E���U��������
��D3��t��HS
]��"�M���2=t�2�a�_���/����f�ꉳK�7[ld���;�ϖ��V_���5iv��Ә��x\��]NW4�c�$J�G4�^N��nl9�
@n�� �oĹ�5u�3�e:�U���=��k��w�B�2[���UnT��UpL�[���6��,�H署o檽��3N�ܠv��$���b�
��"т�9E�Gi�f�:��x��,$+�F�mk�Ҿ��WB=%�s����(x����[Ps������F�.3W���u������A͛i`�-S��4v���ȯ�V�ꡕh�"ٵ��F59�����]Xz�=W���VT�z�qxT�$�> ���^��7�v�\�bgU/��I�p?=�"��ʛ_r��n>8�$`�l����ez��O����?�&AH�7���0��vg��k(�j((G�U
H��+>bA �VP �9�}����f������u#I<�	��g@gdt�gH�ONO�;i"�M�B44�E�*��q�[YXH����f �<?*8_���0~���-@>
g�)R=��:���}(���	 -k��'b(W�P��WӨ3�ݘ��*bO�O�]�J���U3~�@åm>�����i)��.x$}մ79�x,��b�|G\m~���=D��y��UW ��1�����3̑���(���S�L�����
�R��QK�p���G%.:�5��	������B[��̤*�w���[��u<?��1�Vc��1��';�K�4B��YLYÑ��7���p�Fr,�]�	���[+��*0��ԫ��頼BH�z�쨪+pS�)���O��Jz�s!̓}He@�TTUA��޷��b�8/��w���p�MN )7��(���b��xu���zg�:��[�]��b;��E�#����遡�����m:Z���xǌ;Wj�T�s�g_�"!Y�����	�p[�Nގ��e�<�Z���kk���\ ��њ,�H`i��E;+��*...MƍZ��sl2n�'��~}?[G�;�G�Ri�?ފ;�*0s���������<%��,W��4�Y�Z�-x<�ŵl� �UmwrF����2ט�{���y�20PH3YJ��d��)9��7�B""�>�W�,à�>�?-4�+��d���W�>��x�.��u�W�Ѳɮ`��fc��4j�����%�4�;����N���(��Fff
\��&h�&����*@~�T���h'�%����o�bl�2dݩB�y?���͚Jd������&�8��s���^eR��j~��Ū�*V�Ek4��2��٣�`����,PV1. (��k���R�����Fp��ڿ.3�$Au�]�iK�<���w�<,A��U���Q��"����_�����5@R�p�3A��z�a.B�x�ݹ:'G�x}�a��mzͺ�F�ko����Q���M?��@�%����N���d a�j'�pIL�w��B�H=a�X5i�'}��`L��w�h����5�t=6�z��{��B��+1aS��
2������ō�n�~���|ౖ��F�A��]��{1)�}�+y��55jyyy h�V@���{�����WPw��a�Ǻ�g�������v�,�	8�
I�ɊYh�v�{��~�8�\�
��$�PS�Q����{�@��W�޾y�������5"2�2���xu�����(p[�� *u>�|ՖHiT#ΙcC�FE8H�a�����d2fj)N��ܸ���V�;S����%%_��X�A���:�]S��@3ն�����0�ɓ����C�5Pj���ސ���w�sܣ֥���-�_]7M^��z�3�R���ۙ3�-��]�ܪ�A-��L6���מl���+� W��ӫ:��#��><�@�"�����w�eM�fLh��5�� 4�/	5�]����$�W���d!_889}����奤�@ǣE�=;^ǜĸ�9Rj�_��:�?�9	ss�h;�Zb��]�}[����G���������i�{C*P�����2�MK0-���Gg���ʦG�}Y	�0���[�j��ϔw�T��0i�S]̤��(� ����m��b�5?/`�M��98�'�-��3w4��G��, s�mK;;�<Woӕ	��7y"��Gם.G����ʒu��PZ�%�(�7�fD:ChK�0�����������Q�nګ!����߿���Y2���剛ן�m &&4Hح�E����#�*d�qQ��f�Sv�@2f���RN���A:��Z��˩xy5��.�M��XQ\6��P��Oh���{�����q��+�s���v�v�J�͠{���q�"��J0� $����9::����i��fP���D���dZ���Z���z��#�ZE���U��+d{���b-�r�0�C�1����r�>K�{�P/Z��Z��� �N�L[
���+��ؙ��j܄�1bz}yy�W�nw"�:o���o�#_�*a�<mM,v��@*�@���[�gK�K��T�`7�Rj!ϖ̯���Ԓ��e�����ި���L3=}�a�#�t��Q�Rg����5�U{����MH-�ġ�okEn���&X�%�e!�������ْ�ВF�2�Qt�Q�	�"D��)��hB^�t�3ri>�G0�dXx���>/E��[��/���!�#bI����**�+��\�D5e��d����،��b��I�Y��2�kU+`-�rO��W:9����k3���Y_�u�zWY�XW�SD��;�{�x2%����V^q�r�7��#�(pqp2�r�q���J��,���-@����AsQ��-�fލݽ�,���os=�"��H�ϰoEv����xS:�ϴu���N��Z�#�s�	]��OQڀ���"Q�-�c�I�ÓӺ0w����o@
-$:�/����g@�����]��?�����T�}[�[b���ʶXy���F`Y1K*f2O�E?{���?%�g�BXׂ���%���h������v��q�r�>�TC�W����z���Ԁ���JM�:0s�d��f�n`�s�ׄT�d�LLֆQ��1,��h0���ɕ��N�����8�� ��7Z8��͑IC�n4d�����ȗd	:�|�C7�,q�g�Tp8e����"  @CC���]�g�.cl�H�$��p1�<�m�Ɋo��W��Y;���P&m�[��><���.��:#E�U#^��H�k��-�'� ��b��VO�Ji�Ւ/-��r��l�:l8���f��iV�o!*þL{\\���-(�.����a����Q��ꥆ��%�=L74� ��q$��
~�t�y��蹜蟂�1�9�����T�SU?�W4k��%"4?�4O�.0�+3��c����~���i��&�l��i�P^.~G���!��~0��Dfo�7�'WUqd�^%�׿7�E���
���A�g��֣*A�%����h:��^�Z��0J�uI�!j̬<\�Ack�U˚�et��z蓌1b�EP S<��z(��X:���r"h��ړG���r�����j�V�wxH���[���xw�v���D����V| R<�`K�4��^^\�� \5i'��-�׽��3��vE��t�d���dε
>I���+<N���k�Y4����VH�E�O�c�!����Zr�{��RM��h]vvv��"���D��+(D�h�}t��ԣ��� ��hn�����Փ\]���sJCMF{R�KWƣ�vFp/8>T{\ٻ�<h˜o���%P��:z͚x�%�r��=�v�N����H6?�a ����4e~:T�? [}j��pّb�����}�O����e�*���n��7��?y{��hX���i[�YmYʕ�*�2-�''!x�z����vo�֞�sqY�$I�$�?���YZL�RTi��׏��~̤�qB�����n�����$Y���uԋ�m�F㎖��{�*��ü�	L��*�?+� 77w�w"],����,@�g:^M��R�������|0W�F��t���Y��*�%#��#."St�ۃ������:S��K���\8�����5�������k��67<g��pm:�rǓ��Z8::��o�X�h �h��T��T���ռP���c�ex�}_������H�����wnh]]��� -���P%DOO_d�*��BD��X�� P`>�|��� �=��B���wFaZ��n����_�Z#S��J�_��ț��5������{���خ��f�^^^4tt��=iO���3:���D	�j

�fgiU�zu�4j��2* �8~t��"A��L��Zہ�����~�l��K\�V( ��i�b�}��c���`Fȅ��R��q��G��v�f��og�/B�Y�Ӿ�w���\e��F���`V���Ȓ����s�[\J�im��b�(���礥�SPP���������@7� ui:J��/egW��f]ee�ȏ3f�`��n�������Y[Q�ӝ"-� Vm���`r��<�˥u�PhvN�M�퇙YY��l:��bҗ,�a�?�DU��L�ǟ	�T~� �5O�T��n� �)��:�w=��٭`����֥�-b�l�|�}��)quyaa_++���U,h|�o_�v ��&��40<|���/��)sh�z�����E�?M���Cj7G�Q��ja[��ܙ�^ǏH����ŝ�p{��tS�hqq����?0ǝ�@���e#a��%6�|u1˫$�n���k+B������DO���q}��x�uK�4��6"�ێ�Pו�c�>~�<>� �?ߙ ���ܿ�	�ד��5kS�J���rҢ�������Y�^���;�E�2�'���֭����Q�q5���/�v�`wy��ĄX#���/���2�����2�V)Ě���/����¤�:_��#^�7Ş�6+����:�g���ǆ5_��z��"HX�i�|O�����n\�_Y�}��g�f^�-��B1�7���v�%��H7��|r�yLY����&_7��l��}v�*,���#K{�WZZjğJ�s% e��ֳ�d��w�7�����7��YlO�e��X"��E�䭭.�eg����	X>��n�Ꞅ�ǧ���~�ғ922��ݞ�g~��ʐz�?��Y�#CI�X��1��������p��&���׀>{_m"Q����^�-(f��	L+�v�7�J�}!ȼFFF���+��]����	������4?WII��y�3�rw�Y�ةli��LDO/鼿e��""��z��ٞ���r���� FB�$��n{6>�=t�r��ü����L�8ρ���Cۋ�	g-
m�r�Ȃ��$ ݄C�.�{q~��@�4:�a�DbX�,������C�	���IÅ:>f5��>�פ���a{�^t��r$�	�7�o��E��	�.˯�����p9��>��,X���$|W!_-�hT��oSi-���˿s
���3�烼F�+�b�˫�j!�>�-�HY�WU&?~�|��Z.�Kc�,��>��pXH��������24�F��X�RI�sI<�U��Ŝ��B}�:�����\{��j1p�W��4(���&����uj��͔�� 5����Y�E�&�4{:�pҹ^�Eȥ�)(�OY�_��Ž45�����o�r��B�v��a������!�u��1[M���:����?�q�=�Ӭ���uc)�##"��!�� ��A2'� �~��rJJ���xtJ�ޙ���0O�=j��%���f%)x'!�u�U礁R��j��Gm�(�(f��5�4+a9�o!�CM�B�����{�G�(��k�����9 R%M޿O��w1����[[[%�K2��Ur��nt@@V�D-{���ή�r�q7S�� �[F��ƻ�1j�Fook���LJK�l��Y8(^�-�������d��fN�ن��YT����"vA���q�n��v�/��q���cP��\HI!s9,#*�QMmX9�յ�L-�6Z�{���,����'@��տ���)GR41�)(�[��ܑ&�ֹA8 �I����`����e3e]���R��v'*Ǥ��$����R�
m�;���```@�P����/���%��t�õ�J�B������C�
mN�R?��q(��G�pyih�8P�_ժ��S.d���8-y	va=jC�cBӄ�S e�����S�А7�;p��&" ۃ����w�p:W����3���I���8�c��hH�������Ud��w4�o
��v������yA^�}�Uo��>8:9A���/��	c[�ݟ�%	�j%��z@^qs��*���Bӑ�_"6u��� �j���V	��p�J�`�E x�c����������5?\Ǎ����3L�Ra˟��m���\B�מ��� bW)�����"��$j�9��C�����Ы�������tUʳ���F�
���TJ�?sV���TJ�Q�%�`�U����� �wJ9ͺ��4��
d��L �p,=�V�'�$P�p��"�@��HK�u��܃��0>�O$��bqz��W-j��)����{��t�t�_��YG9�՝�����/r�I98T�/M5z��(7U-T�1�>(6!ДDp���Ǫ˷���Eڵ�3�P�A��c��?݆���iYHH_zS7.�rK����c+F'%o����\{����vM*��m'�6�+3?~�Ḵ��|�.�G�1���-7x As���l�^��]Q����;h�-�Ɖk= ��`�L�o�--�UK���Pr�fWw=����5�gU�=�4��#��f��p��r����Q6jI�����!݊~颢�ۇ�	OH�S�h_���N�r�I@j0R��?ȧ�w��/I�x6ٮ����-��g�ߦ�@��1I6��*���,oo:�ܺyq4)�Ҹ�� �:@��L]�z�X{0�/�r�bL ]��'~�� ��5fS�[B�x��t��`KZ�l�el����I4�S���(Y���[���*BB-��B�B�	U�9h��������7���8�I~d���15Ed��jh$�Vl���Ffȏk�yE��[��3��(7�tx��Δ��	1$gv�ڻ��� a645�wq����-�[�P�l�u\���y)��؛�p�ފ�n�d���0(�v��	*��X/ I�j`8 ���Ը�yÀ�𸱻��UP 	�Uf����o�R">��Йgna!'3SH@@`˞#�ĺ/]<lr}h�ɧ�n��F��8��qzW͢������^E�6Ə������bl����M����Ms�7`Y���/��!hg�S*|[m�nˁ!���D�[ng�DF*��+-i��e���y�p�e�8��k=���5K����P����(6����Ձ[�@��2�$��O` �0්���~���4,XT�m:����@�cc\Fn��
�I�g���MC}��5�飴�:���;48�����ᷫ����{0�{$�B������	�xIl-~��Ƃ��	<���hg5����j�U�M�I��瀯mE�綷�w�����A�U��v��9Z���]^]�377��~|_
<�� ��̟�x;��w2T����SV�Цk��H�:�o���y��-ؑg���ْF�ϓ�����=�Z��jU�E���qza@�C�sP�bh��<�9G!/������|�ɒI��>��R|a�/�ƿeI��$���(y?V�� �ѝ���3���P	��#III���sVByQQ(l?.H�x���4���8B~@�x&���'�Y��<��)g6�bJ���3����]�����l���޽���-""x��v}"π�&
���i� 1R*���#5�x5�?t��b�p��<��MIh�t���n&%���Nh�kpp���k /XY 5䰘r��eβO��xps��l.{�^M��l�* a��� ����؆�`*	�6���]�����»)��I��hwe���0��a�N] ��`*�Enx~v�Rn��tq�kZܧO7q���Y}��9�B�- %����
'��"hց����kPA׬�9 ���{��GG%n箦�u�@�Ά���-���g@��K/gl�Cgl%FaW=�Re�\���q��[��)�|�Ғ7�Mn?Lk6[W]ҫb�iW��; �H$n����7����&=׹#������)���AR�J�RQ�d`UO��r��$�|v�V�o�l4a7܇YoL�i��첮��e�������t� (R������<����h�	���}��%�����N$B��'�ru��L~�q�~�W����^M�g-�H���p�32:
0����X��l;Ɏ��6��V�䝡��\����0�a���y���
*%�����J��I:�
듅 �T��`�ѳ~'Gǝi�GP��g=$�iDq��d>�����I@�w%��Ot��H�8r��<�ċ_e���p�g��̨�u��on�y�L�=mA{]���8�bG|e0o��b�[B�,_�O 1��6��i	uA==��溔):k� �AG_��w��v�e���fgcc�Й0R�Vӣ��#:8��Uez{ߡxЉW�á2�V�w��%ҢU���|ȡ`))z>]�p��G�g}��nb$�{��3�.,X�6:xN��$f�i�xe���]�n,����͖G��P�l��zuQ�:25�R��)�����Eg�����`����������X���ǽ4�^1�1d�z�L��,������+��f�#�0�2S`{jZZ����(�-���3�r<��_��"r�邱n�S�5E9�Őw��K�"I@.J� ��bj+Sp/��:04Tъ��ϰ�72*D���2kW�'�ګ4�zy���V/��ٹ�^ׯ� 409�軄���mO��E=G,.vC�j41K\�2b��+������>���T���P}���%Q,Y
b�R��Ԕ�����cPSȶdX��c�o�Ru3�b?άB��'UIߥ��p�w�˶F�}!�2^>\�Eh����Y9�<	 _������ͣc��BN/>��سW17�����srrv��pȘ�+���)&<z���c��6n����
�����QXA`@A`W	i�	EB�;T�:TXBPR�s�!D��a:��� ~�g�����}�=�\+��k�G@�Y���u��Nn9�]s�yGA�2�vonA���|��rF(���}�!��'l�rm�B&��+f�2 E�{q��&��ۋ~Mj�o˺?WX�@7��q3��V�� ����������Vj���@��
b�c��+<@-�m�Ėp�N4H�y*T�.d|6���
V:���nn+_H�\��q���\*;�E�C��w���?5c*���� ��ǧM+|@@ �/y-���M�Ha��"�;��	;�v��o� bf3�!�/�v
�liyB+�k�cU � %�4��q�S������5$$$;�#���k����?䈖|	��q��y���Þ T�7�	���r[��$lb�S6��5�.y�t��1���D �M����9tV��osW�w�.w.{=�(٢�_��@k�[�B���q*��x|tJMC���Bm���ZF�V��#�k	2�3����XĹ/He�t�(9C~Z��i>����� ���x����� �iB�e��$�����\�q���+��sN���{?�%+��)�_b�ٸkW���j:/�+(��!K�ń>�=��%6��0���a��&��~��Ϝڿ�� � ��۫����'��?� 1Z�*���I
?�؏��(ԭ�.�p	~~��z8���S�:�Uq]���^���G��+�S��ώ��&�WhY��=~��rs)�����u��hu�+�s-`'�.h"�%��W�T
��E�F�N��OGЉB��I��$e��П�$��dU��ma�%���@��͸�{M2��CPm�[M��){g�h�i��W��Q��@�:.qtT��TL���=vJ�_)�k.w/#d�s��Ma?	b�Y�dr`|�-��%q@�@9��kf�h����o�=�g:\�Z����Q����]ETW=ڔ����㺘%%��珃]o���|�<+/�����eQz��㛞~�ƃH�˵��<�Q	�ѷ�Ԟ9�-�U�='&��9� |�@՟ W����p�E�=�vhv�Tj,�ݏ�'dA���A_�S�c��Rt���g�UH�I��e�fݔ�h4�ȿ��@"
�B�+1��_�I],Fh�bq����
������zßI�HC�!��.ۋ�c��\��YH�ɵ�R� �#n������[���&C;�����mAپ#1��ֲ�k@fj+ЍѤ\�c3�V  Y�5��;���;� %�\~e�U�[�x��Y	(�����}y{�ѫ���n�[��9� R�l��FF�ம�a%F�z��3���sF�<׫,���
�(����+-��/Ҏ�|�/Kc_ov;��ڛpӧ��|`��h3E#^�ͤ��\��_��m��azt���.]2���t缴�mj��x^��QHL��(}q�UD��x�ɳe��(�yG�޾��N���_!���$0 nO~��ް.U���� m��/]��q���Ȭ����Xf�X�,�Zl�[		�\����>��S��Ijkkc����N%��������K{�(i�2_��x��ˮ���Ίt��u���|Hq,M�.Ӛ�9������� *xK䤜S�)Ub7V���a3�D�A��X����˨ͫ׷��ѝQ�ݓ���J@6�AOx&˿�#Mf�9!��yu��-��E󮯭�9��(����~	6\�k�'ٗ"� ���fs��V�8�t����l������<ɻ�CVj%SXQQQ3����|'�ml5<t�_��N|��YZO���������-��kЊtY��jeffR���\�J�h�W��̭K_`�\m���Ye�� �0 X���h��B�~�����\�r*�W�QW�܎'I����}��m���'�vdm�f(����J� lY ���j4�k���Bh��\�|>F�K���v�*��W�Dڗ`��5W�{�����ņ�"�����;{{qU�_����W��h��+3E���%tW�Tb1���k��#������_.���A~�����z}��io�y]N�OV2z+V�%�M�,�9�sM���A 
�� 	�~�֠8�6---N��Vkv�X�p	�s�K��U�$��⻯�6�.e N�����"%%-��.����T������\vz�!� h�Qh{��k�ϵ�˲y���� ��jۜ����u�������*�""����Ȏo^,8!��1r����5W��U�6 [Z��������Kz6QB6n+ ��#��ҫ6w(_��G���t5�7X-_��PWW7K�N;Z�&��>�>�\ᙙC�M��p��D�����-��i:�}�����k׮up_+2D�,?����c��D�hlUdd���Oz���*�@��U-�A}�SL�/$�멧�G�&���J9��ը�����mY��|e��쬠�b�< _�F����o�g����7���'�m���҅�O27�j�xԩ��>�U�X 6g��U���t=�-' P��ҫ:��.�~���U�΢,��������..���{��/���N�^�_@ @������<|iܘ�s����0�TĀ3̎��/�|�{-��w�Հ���XŚ��ug��nL0�j�/:���h|7"���ٝ�:θ������T؛.a7|��*�^jD��of"{�h��O����VV� �궯A��?������3Dw��(�R񸸸䥧��8��kP�?�7C=9����~
��: �u���|�-��}�A�e�!�<��0�� ����:Sⵉے�r�ܧ.����rv����{�����sN���[�l�G�tc��c����'��
Pe�jM<�ʣ��R�i��6]�}h�"m��T1
m�d�;�������L����}���tͫ)��.=�~2���) �k���Jn=�/(�K	-���o�Tf5��,�S&��a|~˻�B�7%C�4Í�P.5p��&$�g��UX}||��
�Dv.���C��===�8e�J)�P������f��Ѥ�b�ԍ
�q��_D��əW��m�����ӥ`������,3�'�Xb��9K\�I�����M=�A^����}�<�c��� �C�\zE�����Xj����=|����?K��
C�B�/��3Z����x�V� �%�����h�P5���ik�4+�2@@-��X��;!l�#���#?~���h�?`YF�����L��xN/Z.j�[�W��rF�ŭ�|nx�^R:m�,�U:s��̘�Xx=�����Gx�w�������u���bK=���/�m�T��8NC57����1>ᮁ��eu��\���>���>�ap�tw܁�,Tx|�\�¾}u��P��u444������`D[��;��t��C�;k��Ĭ�i.ĥ��-���@��l����g��Қv�#a�%~P��}%��>�NQ���o�'�O�p}mL�̶ۘ*r������u���PϬ��$��mƞ��� co__AnnЯp~(��{�6ŏ�Z܁�(e�$c��g���;p����b�0��@ 	խ�g]N%����i-[K��ד{ע��Mx��mu1��]���"+�"��O��:�<V��"�R%��yg�EJyUs���yd�t�ߜ��x�ĺ	q���kM�L4��[�STȳ{Z2����Rq�&+Az��������e�~.{��� �t?��ث������]o�
��,�Ғ�D�/@�b�W�ӟ��l��~E�C5[��c,�������F����ކ��������{�m��
x��M��e�k][�Y
L��rG�����w�~�1�X���8���<�~�XSǍQ4-�BlO���N�!H<�f7n2��X>1!�+����C��	�6���������* �%�iR� ���xyy��=(?j|���.�N9��g)��bn��?�A�dr�M|��n$�8� ¡��Zx�[Zק���]����C=�Xm@�L�
�g��t!�J��e�_���y���3I�� #,�
@@-3�����Q�ە9���bb���,�5�i���M28/���Tm�=通����&��<��pjq1��H�J��UXZʝ�����p���~s@3E:w���n\��C�߽3�Ϡ�D�vܾ�C�x���A!�ӆ��Dy��Z���l������l�ΝV��;`9Y{V�D��
�	�FZ��yb�h�{��4�(���M�~�����)@ 䓓��ի�� ��6M����	���O����j�?~|

���
 rc3��S r�B���1%h��{{�r��>���z����F2�w튑��@��$�|�q�������4&�SC�V��l�p<��ؾ��Rf|�Z���9�eu�b���d�~y���P��`�A3ʹч� �M+b ������D��y��U�ۏ���koEў��Be�y1�����=�Z���@���(�GXT�ֻ<_�K���$����S�
��b}����P������)���N�f{�s��
����6�-�V�	�{�`R�X�3���Կ*��s��i�'�r�T�a���W�u��j����s��RTVnn�H׸���s�j?����tܦˤ�'��9Щ3�.iz�ȓ���R��K��W�=���t�;r�A�΀�؜��5yd��w���9e�'�$��,�������r���ӭX'�T6����W�K�~�մ⹁)��m�MFG���"�{	�c��!��/�	����|�_�,lY�u�Pf�+j+E��ת�G؍il2YGCmB&6I��뉩1 ��f�bs�G2�	��Ƭ�E����TU<���^ ��kL[��w�CO�<	hȮ�r����p��@%��5$����Pg&�R�R��Ï�L5pGM�>X\Q�l��cW�k~���9�-Z.{xd�"�|��
L�`� JB�E755�ހ�nUp�s��D�L��I��zL�h�q�~ )���E�?@��	�
�ק�0���/0����Ⱦ��a���\S��Ʉщ��Z_�|�R��^�g+���a���o����mf���q\�Ts����������t|Fcͪ�55��FC���G�Xo��(yJ �1���IɃɳ��~'a���������	��p�M�r�` ��E�T%������,�gE'ם����
�@�p}ڴ����g��-��d:|m�'{	F⟧�jj��vZ���45}D���2y*��G*N��HFF�Y�%�d0҂���ϗ��m�lVE6�I��<���A���#����~LC��ag ?�mG3@̳����7cK����&�J�G!Ղ6�RdVJ�͟��-�7F�,��J���r��ϊ���������\���4��K���Ю>>���;+�V=)��B�bC$�0
�������)`�Y[���T�*b~;�;�ד*����o�#��A jU��˿�h��E`c�y��݃����\���rp(Yu��3�{�4�@� ���o�P߹S7��~?:��v98��"�������;	h��?�ʎ�؛= ɺ���i?���:�S�V�_�����b���\MP�X�ho���	��ӜS�� ����wG0r�sPx��~J�����+i�Ny�C������A�{��6���m�@WAe��So�n]#d�P�Kp�t6zx��>��R���J�y��H,�{Ǟ�d&�9�Q��hM|[�p�ЧBwsZha*�mmm����r���R#.v�sѧ��T�0�� ��ŮM�e��Z���]�J�~NuI��������&'��O�]#�b���eu�GZ���K/� ���f.��چ1�V�t��%�����#�q���>.����#i�V� R�K�~zP�t�Bsj���Qs�ՙ�D����gb�zz+-	q t8��<c������%당����_�jr7�O��
�ܘ��m6�t���0�"�� �g4�!DeƉo���u�������%��m�;�iil�>^`ޚ_��C�0IZ�u!��ֶ��6�뾚�.��U�k�BJq�	�,	�����>jض�F� �Mջ,�SMZ��K"ƃ?��U�"Ϊ���f=�Feo�]� o�T,ܱ����8�|�|�s�s �l�nE�;���=��-㍫P�����4}���V����!�N�ZG�CϪ�)��q�A=tWo����0)5F�j��^�k�/�N��A��6|y?�}��.���]3g+��I!��G� ���d߄��& 2�d�/���}���3<5�Nq�=Q%Xw7�8�ٛ�w�և���O��6�
��04���oBB��	hiE:��_Q��ʑ�W�Dj&=�W�%���q�2���ߡD�9G!9�2B7�D1#EW(���~�� #2T�o�	܅�
���M9��!򖆏���I@^�S�ݏJ�Ee��M2��7DT��A3���հ���P�/q �`�����to�\7���:r�aKDUom-�tM��rk�̖��:L%����
 ���'��'rF��/���u��Gwɤ�]7l���zyii��A:& �ol|\^ ���}[������/��PNz�'�<@	�p��/���]�:C	p �c��GCn6����~�v���xI//��|e9`��A�P�j�q�Q�R� �����%6�s��gz���\>�txP>'��	D�4yy���cW`*���ꛞ�w.�oI��TP�=���h��Z�D�tYHA �J���*_��Y����#j��'M�->c����m���V�����G��H��Zh5ED
z��м��˽����e�e��ֻ�%�$�2����2W��&3J�CɇP�E2Z�,��TBR��uIWO��S<�������ff���wP+���ܷ��&�����s�,�����2y��w-�x���W� �]�q߆���jƋ�5y#;����o��X�_&$$,����0��o��jV�ag��@��5�[�
��><q�D6"5�$S[ .�ᭂz&�T��o'l3~���$���R.�����XĽ	�T(S�?�j���'��!"��>����~���:9�'��о�u~�*��[������]k0➜��{B���
9J�"ǫ�����Z�����.�w��+j?0�ΰ��o�@P��|VΠ)��p�ky���r��wtxSխWW��]���X���r�mm	@�QA)��Gc�J�#W{���~ǸC��&��'n�8�����U�8����-�"r-�{��׾��&��៖�gҬ���r�nvY�����';h�=�GYZ��Ą5�D��$ "	Ll�J�����E�
b\^�:�n:������Q��笢���=��N�i��33��z�>�ی,����,)w���2Be���;�_���@�^s]���dӿ��W�t	or�%��C=�(���q[��蟩p�o�C�lBb���Xf�%(*(@�����m)	h2� Iy������l+�"�گj.O���ꏡ��S��/<�S^ {�l�U�p��i9�^;a�#����I�����*���F	 -��1���;y�c�Q- zɧU2|�5�1����� X�&%%]��G�-{������m4]!����R2<�_���dQ/-�$	����+ ����:89�ػ��� ���ɛUu��h���2ޛ)x�7��4v�C��������!�?ۡ��3��v+���\wu@��N7"V�|��Q(�u\OR�t�IB��Yf��0�"��?��$P `�Ag�7Jo����I(���B��V/�	%����>R����E�6Q?#n��T)�o����|��1Ҷ(��6���*�sobW	�c�*�^�ܣ�3���e�<'p���aM?����bW^l���#���3�S�7�{M�ԏ��݉~{U�Pϕ�V��n�0G�ޞ��C০�{����:���5�`�K�Fj�>�])�n5��p8��/������%6�* -w֣���,DS�x�+.�G��E�w M�W��e�MJ��Q���.�(�E��w��ם��!�����-�����	hy���l�;n'�_`nN��ןN�6(���GD�<�K("j�_ ����W�;�ƅ���7�|u��u�5W*d�VπTw-1&S�p5�P���ӣ�Z%0�>e֓�?���ho]�+ ���/��AOJJJd� v�8�D�JN+��[Xu����9[U7'�g�.��&܀'�h(��_��|r�б8m'p�T��=s��,=/�M�<>@m,i9e-�l�F��ĥj�`���Z�;�]���dVc�L	��W���H���C�\��˳�#'��s��y=�+zQ�zg��\�/	�f�s!�}8�o���Z�Ǧ��<]�u7S�s_��'���O.���եde̬sv��eX?��/OZ[閨�ϴUWd��8SD����(�Y9W�ڡ�h�����
�8�\s��Qy�����dd^^�pZX�hyOr2m�.n��}�Qv{�Y�X�ʆ	��o���h�r��:����_%hԕ*On:�X��I��^���+B���8�Z߂��ƴ�J΂�u&aq��s�!��z�(���^���4����\:P�R���W>��y�/��6j�ebbR>�f��Ps~�Tj9�~5��(:�N�����ӡ菟b?~�Z޼��D�Ip��bi�N�"$��߼�l�s[h����>������TP���[�b�4]���X̄�ƠG��vla_զ��y߇�'4.E���?���m��.��ژ����*�z�N�(�����c&Q�l��9�:Z��&KT~T��1�u�f��|c���P
�-�������+�=vJ��c,���dTT���	<�cy�W�R^���yj�0^b&¥3դ���\��p�YpEPh�q�6�NQz���*���&�#>11{xV�CQQ�������On��#,L��������"���´���|[r)���������=Wk��s�|�䭭�X��Ӡ��96ぶ�4���~���s����)���1t����Q�t袰�>>��呷�/�/{>�B���s\8��gs؏gR�3m7,�)�F�\��?���i=�5X� �3� ���Ne:
�/�m�Th�4���fN�	����E �/h�nz�{^�7��߿_?�!<����ޥ<j�}����NY�'C��������<Z7��>A��yz+D]����9
������";B�~M�Q>�G-�5��R"��W��7AǦ!����<��}�,��g|��'|�V3���o�i��n_o$~��5��"����ji�ٸI7g���_� W3�`~ۙ��?��B/���Y ��a|�XW�݊T�3��<C@�R�s+mGyD�V+���s��;'#�����{��/����˨F�\RRצv��h�Ǿf�--,�`n�`fR3>�2����A�+47*���՗��Y�L���j�N�,���{A\/������b��}��Z
�&�u�� �ֵ�����1G*)+#���L��X����}<�Urn�͈p�pu,�sy�VXdW�L�p���&�����t/Ĉ<��!�W�41��h�z�tX����	i'i&R��Y����h�>O$n��)ؕ��[3�jg!*��د�/�@�w�G���7�.8���	'U��ї�46��7K~�[��.����ؐeP�f���	����(U׬;����潴����}����4�'<%ic����/R|��K�[�/��2�4�%������t�?�-���֠v��2��ٵ��Ղ�C�yg����Y6l�#خP>��yT���V4�k�y�4g&$5G1��ѷ����d�E��a:� ��?�Xo.�8���9�M�z�D���e��NP�Q���W(�0'>.��į�SJ揮/=91�/tO�E���#GU�J'� zk�A�}�߸|?jz�����z�1GFFf`ż�{��i\��R��Pl:=@D�����k���/�~5u�N����V�T�;���4�=�/?�3>�.Xj4~�ߌ�"�L����	#v�a,zsb}���9���Q�e�JE-���1����u�|_��3�֠����������	�6�$�?I���]��+���|��u{8�����K�T_�(�fM��ҋ2'�d-l*����Χ��WJ���ti���1�<����(jV[G7��m�t����o�(�<��9ڵ�nh�ʏNAn=��ޕA^�Dlu��"�i��F��j�~�3��|ւhKu���(Y	:os�3�5���\؂�$mr~��I��u~N)�ҳ�I=�Z�O�7�R��I)��/���b	�+�M�����xѫ�X�,?����ou���LB��Y ��ݳ<f�8y����L�*�	a�fqY��fh��kUII�'Cǃos���?X��{�"r���\�e��	�sݴ�ŏ[�d2,R<�O�MҒ�������t2F%{'�����Y5Y^\|p��7u�3�鿯rw�� �)�����.�?���,�����DD_�����CR��E��b�w��ق�eZ����Q�Yff&tpxtT�q#�Y�
�M�����s���<�{]�)H�hyK�[=���6�]����y�lyg>��:�|-.<C�%,����t����^��E�I�R���49�,�xd�bO_Bo�e�@Y�@�;J���}^��@�J�i1��^_,F�i���Z�i_c`�Q�`��i�(��參@\k���QZ֩���Li��]�{dx���<ϔ?�%�ޘ�������9�Gd��	b�e�A�s�{���(�NN��{y�(�a~nnGu�g�J�P�����[�)�߆��U����3/MӒ����C�yQ���)0���I�b\˶�*:����KxXB�a%�BJ��NS��V��} �R��j78�(4��`Ek�0���Q��l���{E,�Xv�v�9����[	����u����:~����-�e��V� �5�9G!��:�R�o��l�_OT�:��+����Է?a0�
��b�`���
a�������:�b`Cd�A�L'LQ�E��	9���+Dr��=��[&Vv(i�2�a��rL��6�I�v�}*����V�s���h�S�W��q.�	9
�!�iH�u�wƵ@S6���G"C��#H'�G�U�9\�Z*D�`�:ۯ�z �M��ٝ{�K��RXZ��UzkQt���X�����,�|���K�[��N���cKt���Y��
L��R��A�uO{�k�ʁ����d:O
�9^g��6����0~�}�I��$�����Q��5OvBGQ(I��""'7W�\vF.����xſ��ۡ���&�`��~���~K����?��3�IN^,u�Dz,0��2(�ĩ.if�=��e��F�?.���J:���o��BTkP��}#�lOLa�w�����p�<�	��31''���gW�>��9�4l�6W�PX��_�et�)T]�?.%'P~z�cdd$ݾw��y�s�+��n��6�����Q�9hP3���� �����J��D{ �s�;�A�K���Ax�Ό����{Ή����Z4NCV_귨�%����	���xG[FC�-�����6������"� ��	&�������������U��!��qv~��b�#z�l�����p�n�,;�߹ j40���c�70X}�E��T��vy��+q�t|0��L |�W�/t�� �ݴ�D�20���t��þþ��F������0�#�r��;��F�&��'�����^�]�a��U�H cGb�_�R��]5u��w����#�宓��f�C�|���/��s;�;#���L/?��G������`�/	��8�x�V��%� ���mv~x=�C�$��4bh�b$~�ޜ&Ee��`*���9�B�:�9�^{ˋ��e��V	��&�\(��k�"u'���u~F����꿚/��Ө4w��]�rV����JB��j]F!�����;VW�T݁Հ��!#d���?�����ӢGK�x��l�x�FX�<��i�3�#�yx2pZ�y���P�*p>�w�N5�z>�%CM��GGu���Z���
ݍ}y*��i&*Fw2(�[ֵ95翉{4��\w�w�牊3��z*��ӄ��۔!�$���fuN����ca����lJ����C��+������C�"č*}�Ӏ����������uq��)m�a��/�jg���j]� _����dq;��B�D����J�ˑ�]K�]� ��Bi�D�.�;�����vK��7���>=§��Qc�^�i( 3���5>��1!��m���׏��KU^)B�y�
A�\���.�Q�+���F˳������,Ӏ�`��ո�/_�Q
�J�~�\����Q��]|<`ݯ�a6���3��G��~�$ϔ'_���u	:)�^�Y��x��We<뮾��jE{��>�.���K���5R�Ni�����d/uz�7�=M�'0j6��oE��փ�f�r�؟?K!��`�~�m	OB�N6��/����=���Lu	&�Sz��w	�M�Y+sQ���Q7�b���)��x�$%��<���V\r��po`غ\]���bk�ͱ�Զv6�{�X�ɹF��k��4��t!#�tlw{�enș'/M��JH&@��%o�|�9�1�
�Ha�m򡦦.X�[��8Cgĸ��;�G����4ΘMIB�+��jօ�������te�"�� �ʔj����s e��5C���~�����9h5�x�M�F���>!7T�^��/&�N�e��$�|�q+,��?p8<�__��p�/4Iȁ�82e" �c_����@Y��t@p�$ә2�, ���N�J��YXU�|�4|���B��BÑ�����PV��tr�����,�
�9Q�lY�õ	�6��)���B'f�$�_Pa�4����f��ù�oX�h��[��v��]B�JP� ��"�*CθX}�ꃗ��o��w���٨�^g��B"�6T�;��t>5_���r	 wyΘǿ��%&"0�@�c
k���쫸\~	�<�0���a�'���3����_i�N���o��g�X4(��+�!�YM8���`ζZ?��'YEst���ѕ���9���+�ش��P!���6���EF���H���~M��*�p8tt|��@��^�wh"���tJop�*YN)���4oF��ΰM-���O3�`kF}9B-L:���'BX�5�S2i���}�\L�ŵ���6�2Gկ��}�J��^p�P�A��Q��`�{���*W�v	|��F$v���Ȧ��^���f_��VBk�T-��h�Vq[�0������ ����[z#c@�G�ǽ���d<Vˏ���۷���]G�0�D��*ӎ�/O����:�=sa����%u��(����~:���p�x�
���**�!�
�m��d[��[����'@x�>vW!"���
_�GF;�њ�6��>;w��kw6BP����M^��bXM�p���f��I{8K�KƹW�	9��GvP"`W5��p�p��y�M���+\@=�>a�6����.}�eX���%ӭ���Ac-����/�qo}[�̸�&\zV�Re���f%�k@����^p����E�7��2�M�}�)/B������w��{�>�ӓTh�=�mR��nge&������o������!@��pu'�|�-�w�r"�,6�
���^��{��	{ƨ�/�?[W�*W�*��(�P�:d��?!�� U�p�?��3?*A#$������������5���㓅Z�����]�=l4~�ݔ�/���⮮���ץ��SL��Д����	��<\���%���4Ȩ��`�/v�U��\����~�0���������S���4���W g���eW���G�W���+7ズn.������<�į��-*��rg<_:�:;�L@�����9�`������U:�u�L~�u*N���������x�Q�ή��#^��u}}QΜ�+|��z M�u]w)����9^�� �hɂF
u�G�|||��YlH��P��&֚qßU�UW$���u�=�3�1��h�R����@\{��gʾv��.���D��V���B��W�Q�S]@򟟐�J�G�<��&���6��Fю6 sU� ͣ<�3a�a+ U�E�̴^%%'G��w�h�Y�R�&&&���P� ˂�&���L�uN%�ӳa	��=�=l"^[2�ΣD,ഏ�Kh0��z*.#������DН���8D�Vsue�b���meC<zn��������B }?74�7Л�J}L���1B��H��8tw��o`�V@�����WBэ֛P���v�\�84���#ګ,��*���8R�O�9�{�;P��{��Sl��q���v×�5e#_�(/,"ҭ�fn.��>~� "=�(���X�:5�����4 �)Ӵ�����H��w��nŋ���dʙ��}�E��Jko��Zr	��$ ��Bm�����e��NC.���v��I���ț������W2|��n�,��������%�UPm�< ��K���r�j���[�Yʏ ] �vwיv��,���I���I�i�O�|�j<��^1�Ku�A��.s7�̌�q��$&nT��8R��b9 �	�:;%�vQ��i�o�T#�9
Z!Ǵ�ܲ>��%έ�o<;�����f�8iy�W���ᖂ���T�T�f��+Q�U*�����t�:@�#���W!�Ζ���X;��-����:��hHd���k�3��S��N�ﴂ��*�ȿl
�Z�r�G;����q3��������������o��v>Eu�x7ǚe��}m)��E3�9Ң��ͯ�Q������ps��?6�>PfVJ�������X3nO*а�r�CM�5�zB$,tsk&��'��8����G8���*uh�_ٺ�&����}�6m|�Y߃*tQ�{�Nrv�"�3�!%#���)�I����6�.�,Q�&^�-������̙��Xe���lk��==k	))#����K���m�SD�q���՞omgg�k�No�:�@�˂%e}��->|	��i_Ӎ�С��6��H��о�|$�8M\MA[����x��G��@��E}T�-�Nq �w�3F���<K������)1^��A5='~dA���2o��&��ع$is��<|F$911a��k�B��c�T����!�JHDD��0����d�z�/>��%���$F�k؀�� �+?x�m��ۂ�x}��{�tW���j�C�Ru��/��?�!������x�B@� �����mZF��j�&���S5j�X"����Hڻ�^6Ϻ�������$g����at�i��}�UTF�(� �@��`��]�q;U����B��{�����i����ǖ���{�Q_̣x�߬��>e�*'���΁�ׯ�?���fK�ק�
���GE[f����$������J@'#t��OKLhDj�Ԙ��XxS�ax'R����Bw ��w5hF��=&��ݬ !	��5er�	�H���>�H�2��\�\��	,Oη�9ǁ�+��~�8�DT�T����]N��p�+d-z���P��)�;�GNNN>�4�];�c7��O�������6B�B�|���Ϝ?�bl��L���g֏��R���^9M��Q��I�uKV�o�+	�2����u�����E�U�udј\yg=�Z�k�l���pS����[�l��,��i���_�������Ϙ	Q��
�����<��|�4�S�׏.q/.-��a�I��5�R^�09�	

rX����mf��=����-6.~��:[�GM��n�.dV:���談6^(_�A�7w؛��7��%��V~�P�э|��a\2��M�M�v-�WՖS;{�GM�-	U��0�Ǐ�S��n޼	��kr��>���ܕ�o�����|��nC����q^-�x��?�F B�-��ݰ�.�,dH�+J!-#C�r0鵞o�)R.ho��1��(Ǚ�D��	q���s7/�=X�pf���Y�CE��g_�n������j"w	f�-��|r���,�}wL��O�6.Tn"�|�J��ի��_��Lk/
nŽ�����ucœ���xz� ��tu ��|{5��],���[�SL�Q�,��R��*�z�m���w�E����m
9������O�H@5���� ��&
�K��eX9_� �-
$t�I����]Y��5�MP�
�E=��{�n�8��Y�C�^���ww�e4��bz�'��%�+�`ħv<)���eW����=�g��ym�>)��$����faa�{����Z{���p����.���/vTX�* �m�����ָ�\�M��>'�eJz::y��@�Px���/.��$�>���t1%��k�9X�J�H�Z?�+��^9�{� Z.F�J1^юS�V�������?br��3���b����ZՇX]�GF�BG�᫈Ɗ�e�v=����9S^U��G	�D����1������f$.�L�G��,]LO__n�]&����\,\p0[KYc�����;�k�a�U��egg2[)����w4BK[Z��x�:�\�ة�_9�V&�Wz�� �?e#�ۼ�W�}���dffV�Y�A���1�$�eg ����s������;䷉�)�2>�O������L	)�We��ލ_�~o}z9K*5�2����>%f{���Û�C��C�:�89t�99i�x�j|Β+��
 &��^��s|T�7�sX��ܷtt�䫕,W�,����) l�t�X&S��:f�������>����{3v�5�:* �l; �y�) S�����$ԃ���2�����u����T�j\Y�r>�n8���N`��Gj�K��v����~#?~|R˿u⬣ma�p���8��!�4F' �n��}�T�1.�L+��o�aWLED����Ǯځ�		I�zh������+b��{/b'ȚڟK+�:\�Pܐ߃�B�c\��K�Q0�~�(��a�5f[�IG��2"��knm4�l�K�5&�b_kO���j�ʁGӊzj\@\b�������8B-�����~0����sg�pZ��_߰���IM�
�m��v���"\d��!��2�*Bv����lb'��4���0�[�z�/m���]�q��|S ����MB<�m���+<�w�������ٶ�`��n u��l��ӿ ��!7��q#`�ç-��w��;�g�G'��B�V>ՠ
ɯ]����rB�33�Q�!�]��7���-�{{	).�^ϙ��{�o�q <� �İiC��|��<h�~q��)��]��lx�?���Y��2sD��A�e�Zy4Q��@D�R:���d�z-r��|��̎ҟ:U�(�}��<�>vs3M�p�#/��sKˎ]=�b�2�a�����V������gcu��zU�fvĝ�!��� ��k��Ŝ	���_2�X��[oF�4��e���W�{�5��ƨ�?2���7��dY��K�\�U�?	��WW+�=ob�4�M�� ���N�i�e�g�#��z�U�D�%�2dXO��l4�pl7qSP��j����֭�o�p�R���zR6f_l �ӫ����� ���pO��]�T��8��#�"��j�q�'G�f��+8�u�ʘ�ړF��0aaaK^�J�d��TSid�p���޾���SzZ�M�$�j8����Hz�b�+Ā�x����k�����hxbb��.j5��Ғ�SU�UĿ��`X5��oߤjL �U�}����N�$d��u�aMfM;ꂫ���"��T�w\Q@zG�J/�C��"������^B���C@D�I	�tBB����~�%?�}w�9���}�s��H�UKo&�e�Ϟl�}���l& $T����e�TY��������9�Qd�̯�GTp����(C�\:���Qz�q��\�cy���ّ;����ؼ�����%��	:,|��'��CoK�)��pD�j|�#J���jq�:���[gQ�_\RRQ\www�&����2~E��^]`��!i�����2Gޓ�f���$�g啕�_�̅�ea�����a���_ �XI��]�u.�^V��[�o�QÄn"�I�}��N�1�� 7�Ã��l����nTʲ1�%�j���Y$0z��_#\�cC#��H���eM(M�0����zJX5�w��s�'L��ҏ����4�D0���p�Q��@l'	H���R�ԢJ��o��q�0*+ݒ2�!i�$ͼ���t���/D �Rew�.�+�>(�����'��t?;���\�����E��z��bf�߹�08j3v����� �CxWb\gIH%�{y��N�XD�o_�~�<}�9�{������kc�9p ��N�$�J�sC �4;;`��,��q&{����z�<]䔑����;�����t�E�Y���P�SE��ڽ�ܞƋ���,��O��ݝj%�j��:C 5��p���7�VҠ�L�a�&&S����j�T'n͜{�\�����hZHXg~f��hg{{�����I�f۠^��h�-��`I�LC�s�� n-d߄��T���]pdI�|\��N�&/`���_~<���~o[��ۊ
>|�sV�E�w�τ�uL�?}M�Do��:���D�9�������ꇠ���I�����|
�K`2{��N!�@����;�T:��..�����Md��y"�G>跷�2�ʋ�+볲��%j����c(�1W9���>���������p�����vN��Q�h�����67���0���Oa|#Y߆XܥV�3�4wE?��;�QMoo��^G�pIn�_�*X��;T� ��A7����
� �C��"���3g/.�d�Ũ�� �87��ep�b�&���r�^����/kNtWF������rkRcufZ��c}���[�+�g;⅄�r �Vxs�Hw��P�\7q�o#�jܳ3�V4�F��6sA)��bêvA�*�b#�&V�����e�D�4�"}Sά�_4:F۴s�j�d[ĝ/������>4My}wf���9��4��Ѩ�����c߾D}����xM����Pa��-at@�gyJ�\8G߂��1�o:�v������u��|��/Guս�S�$�aĒ���b��B�ޞ�~�p��p�J���;]]]�׽K�|fq�~�b�Ĭ�D�N=y�~R@��{
�H)%%��� �wG ky�HɌ�õg+9�"?߮�ʂ�˘:DY��#�a*O�Id|v�Ī�q>r�U^�Y}zNEU� /O��<Z����k��p�L*_܇�![�����i�I 	�a�gΎ��4�0 A֛�Q�WI�-qƾ�&��w!�8����5~D�4�*[�NS�)r����z�Ɗm��g�aLӑ4\��;���N+s�� f&&'������G�^jz�.+����mY.dGgu���!��Ë��o@�r���Yn�^�}��_�v��U��$K:C<��nZ7�ҴP�g����\�Ipț����-$h������� ZS�W��oit6�9��4���;X�N��ϷsrR�R�])���\M��a,��c�eQ��9pt��p�k&%w��yڽ��謫���ۜ	5eX�߄cll�r���AqBJ� ԥ$��*D#��?�u	@�(c�I�J��e�����S��q�5�{B	-EA���'��G�l�O�=mH��U��G�K>���a��@`u~�n����\-�k{�o[�4;��fu=?k����l'|7T���Π�����Tϟ�f7���2n��˵0kkP�'��2���&�`��uP|�Sv�a�`��]�3u,�ք�@��\�� ��2t�w-l�lncn���d��4?p�Ls�C��s�!YK�ok�WC~���Csq���g������`f�郌4ws��EX'»L��ߒV�n�C�)XE(�)����e��nU<����n���ɯ�$�-���UiUQ&h@�o<�B�eEmzU��JRB���`	7�N�_;Xa��8˲�#�1X�]��LP��z�/���e�r�I:��Xݗ�qPe(+y5j��-q��]���Ď�Y�d�G���
��56M��}�g�pU��B1t��&M���O��t��e��/0X��\�:�!�"&,-(�8g�j�V '?�u;�����+�1�݁������i(��w��V���u�G�,�+�#������Α��ϑtk���j�)))��46F�cu�ɇ^��݅��1_=�������5_)��p�]���7`���V.���dv�޷�P�(]�}J���IIZ����i6a��. �����*�������a �����������%��ס|,��ϖ�ĄI��������e�>��	�i����ЪR���4|�h��
�ņ�}/�z��@�P���4����!�Xd1`Кyʩ���pY,!h$�����A�w��Vby'�U����g�{L.y�����H"4�%�����ydVV�����-�<��:C(bG,�ߣt��4$R�jj��C�(��Ih*�Χ�����\��bKb;��B\o����q����8�$�p�Mi�Aԋ�Bac=Ϋ9}6�m�7���["��2c�.\\\#�pC"E�6�=)���~����+p��kY�����<��@V���["�uj���R�V̉�x���+.4�vd�-���5��L=n^"B����GFB�� ڌ��54�T����<"�`����⧅z����?��W�SN�<i����Q�xr�D���>E�Gj:��Q��l��ɭ~-�rhI��L����N;�A�ѳ��8}������h�{u�gaN���A`ͳ�J��ޗ�TƵh��i��X�(�#�s�E�-CwP_u\�1�YTz�Mq<����/��n���>A��p̈́�;�++g;�(w��Gி��ϧ}����Bj�Wb�3w�}Ԡ�Y6!����mK��
���1�(:�3��J�b���t��b���3��XIUG�������~lnV���`�wQ�B�if]�h�~/���D�i̴��f��>�Ӌ�`˄
�|Sw2V�����x�Ӗ�F	]}iV�ۿ�X]xS�g/�<˚��nM�
3Bl�`�w	����
5Y}�h�sX��8@��P=��׍�v@ެ	�8,i߾�H�=^s;%����k
�}�Tu!\jw��%���0��u�]g�d���	`9W�w5�NzgQE���Ź�$C���N7��rz�BmH��q'zdS[��i�
����q''i�G9�����<��ı�\.eN�r��X�W�V�.i|Em�#���c�ӵ9��^��)�)��[��V�� �rP*�Ø� _����"��^���lo8(���K�����6�f������/�2|���D~��>�Xw�/�8üߟe�p���=�*�%(-�����궐 �V�,��bF��`�GDK�ߧ�jN�����>��l���åB���1�u���6�6!/ �_�gB	�\�3����źBbbP.?`ٌ Tmh�d�"z�F�3����ln�i����o2��'l����߯=&�ӧ������2(��.
}%L�<��u�a7�n���y��ꆧ$b#X�
�ߚ����<���([�<�+�s�������s��_�h�Tt�D�K����*���*���@�	�6���R���k��O�D����C���J��l��:<\�\e3ۑe�AX��Zf
��93sss�q0N����"�	Y�U����7��i�W)�������0Tj�D  py~�#����G<�ħ��e7�m��{k-�|2l�,�`�Y۴�zTqLk�p�G(�$���4n��3(w�E�5�}��ٚ���q	����MC�0F��Z�ow��A�۴@3��QZ��	d�=�FE]z���v�=w�� �رmB�Y9y���P=_&�j�P�������*s��W%S��R���uwG[�}5J���� �ѣ4� ��v8��� ɺ����\d����Uw����GeJ� �(h����TNS��R��%��Z����A14<�J�ރ�K�>��vZ7�S�}im�g���o�ӣoxE�z(/Dz��#���ɸ�������Z�J���?v"j��(��,�*�<�τ�R�7I�v�1�>:BͩJy�m�.�vԿp��[%���AC�Ž�4=@��_w���X��W�$��ckҀg��c����ts�?�RT�q�lT~?��p*=���w	�x��R�s������e�U'�@�]ϴ��$�"��[#���w^��<�ӀQ*��bXz}��ߍR�⢢��W�N�Q+�b���q`8�}�p.����[" �(��f4L}��\�]��U���M"8 �w��m�֥�:^��k�F7�)�+m�ėo���Ti7K�*2A������~�#9996$�ٿ~��'�P[�s+��;1OS��ۃ[S���f�R���(�����| a���]p0��^�Sк��!���4�cM�Z��Kn����F�x�+�a_��IM������\�?#c��#++�_f�vE�����:���x��ZE��.��J�b��DSW	@영��w�Y�S�u��Dg��r2m��au��������Ss�l����͜��,�М|?��QSV��	G�e��[.��J�+ԓ����A��}1�Y25\�+VxS�07���a)\d\���Y"��.g,T�ݔ ͍�YY\D֙���ct����v��^��x
�,�#���xϱs�OO@����ۖ[��{�5�-;G�����E�i��G�#[�  ���y+�Ń[h ����6glE����z,��N�_%��������퇁>u���-z/3��sgEչ-FC|�eУ�U�顱��@KA��g{ٹHs�t���Q8��61t�6ko$�rZ�3� j\�g�V�Xa�$��@����w��t�w�UǊ�����Tˍ*� D ��}s�]w��r�G�F��Y$�*����0#w4XL���D��.�X_��3�j.��d�lE�{����f�O��hll����-pf�:��H.�fl5��8U�����,sG?N۠fɃ
�(�����ClGױ$�^x���؏-���;���f?��g-�OKJ�r���nm��H���i�[ڜ�vV��ꜱ�2B��F}0޾)����ǁ>I����|��r��ˋ��%N�ܥ��|����VP��1Jl���V2�-� #޵,M��օsk��$��1�)��r*],!������	ɳ��Ϝ9s�2hVF�D�ߑ~Pp��Xe�i��]�ez� ͓�^���xs���� ���pW󕖖�D�KNA�;������g¶���%^�&�?��M������w7E���\��  +ц>*b,"�#��\��Ãj�3�Y��c[.�b�b��?��������v�wĪJ�&K�j��F�'�$��TJf�6���c=��&�kO�.������#�<�Ӛ��������+��n�����.'��O\�������muDĈ���!�5�R q�D"�
}�[�`�~F:Hm��Q��T󶠧�Q�,����WF��c*J\�ۈRk�b��z� #�5��YjM�̃�ڞ������4����I�X7ť�$[l[qҞ����cb�*V��\UĔ/��u���RQ�'�eE�}�����˥�q�Ôp�l���&��G�V�ǲ�v��_|�˭��>5����ig�i��r���@A��6��	*N�k�+O��t��%5k�Pv:���"17..�m��H>��-,���M������9�?��/�병:���e�,�Q	]�I��k'*�,������"�1��/K��	+xLɄ�� �7����m�W��8���^�mm|���������x��P��q��� ]��|iU.���?3����=QNb��&U��H���6�J�Ӂ�3F���xxx;E&��bw�:o�#I��'�o/|�0}�/����NC`��nٛ�D����\�LǸ����'
�1[obTbq�;�{[���΍b����x!\ _�hl�tE�h��:��ٌ�<��P����7�gM�@�2�S�p�Umŉ�]$"�^��ޜ�����l@&+**�	vn�����饥�h6s��~}���?z"�b�4��2{12�7/�|������E�3�=ҳ���B��a�i���w,�(-��7�/����L�`�kz�{x��##KvZ���da鋬<<t�>���ަן��h�.-@�:�~*�ʺ�o}�D����*�rz�k�}{�y��S�*b�"��HU��I��W���I�*��K�p�ƀ	���n���_hg J�仨I�}*�#�����4ռض�m���⼴����
��ws�r��5��d2�� �۬�?�c�ҕ.��L�X�)I��&�:>^��&��}+j�vd�L����Alŭܖc=NWFO�#;��	 r�q+k�0�^E���2��G��񟐜�����X���l�;��κ�4������W�|��'����lB�#���.��1-wH�Mէo�˄<Ѐ�N��!`�W��NU�m���%�F/[&�BA���m��Qk Y�>�彄���HV���k��(+`��-��3"�������`K]P$��Ь����D�ؑ��10���iZ��j�">@L�&�J.�����C#��{����;��ڼ|�yP*���{����"�	��%�Xׇ�!�e��)���k����*���أm�~��������V��D��Ϭ�N5C��wv��3L1K�_��x�{UW��S�ȸg ������5�?��ɘ����#��\�z��-�I����=�@jA�����É%;L�������)UI1|K�����}�9C`�~&%(�0�.�
�ٚd�ܚ�)Y
T��~��0�"^a�>�XŜ��@�%�>Q"�J�B��DL��ԙF����|$���P�Z@���76������)��N��&��	n�Q~*��￙�j�����|�)�Չ^i����:3YenJ��twFv��8C������r�`���`#A�u��#��/��J6��A==!A�l�Cx-���\�i�[0� ֥�hv�j�'��x��ㅟj�>�9�rb#�&'���Kd���K�=��O%[�A�Е6�5V�͡&��Z4$�i�ո�l�ގ�+W��-\sDq�}�u�p�0��V	�co�Yvs��m��5�%ٸ���I��0r�D�?�����b�9���Y�� ��bccC�u�w�˷�������TF2��1m����B����ݐ��{4�ׅ��">�H��p��N{{{붡ܯa"�L%⬼��k�J,����~�1$����^Q���WӏQ?Oq��n1��'IڷI��o��v{ۧ>�h����鵒ޠ'��E+A�#}$���o�����߈����:}pC�}ˉKVە��9-�裴9�'}�1	>?l��V��H�YHٰ��1�S@`fo�}�pQ\|<�䀔�hl�TxE��;}x(;�B�O$��L�%�?6�P__Lʓvbz~���H��	��0�%�j�.���`��7��G���1�|�����"��$���)����1�b��������9�s	�o
�
��k��?�Eyy�!��J�|���ٟEl�r^����x�sd,�n�(ieeu��;s��yI�T�⦪��>�۾5q����j�$����_)�R��bMդ�>�\��;��9^N�Dz�2;�[�:~:��}�����&  ��|6j��{�5|��>�dlYq�4���_%�Oݕ�Bg�o��́�S`�<K�D�m̻O}����jxX_�36�.��o��q>1)�=yO�S{��4��I��SZ�*��)@)wJ�rfOn]�;�g������)ԁ�q<���@K�$~�O���?M���|D�0R>�!?5	��Q�%j����Zg��{��<�\�[P#jq�-amN���U���56�?%F5/}�( l�я=����D��	���`o{n_��0J�s�|熹�IZZZ��,J1'3�b"�������� Q��r��g�K�Q�~�RLO�TW��)K�z��&\��@o\����U9�|6�+�V����ݲ��d` ̊�(< w�D�W��t�G��]Z#
#���ЃT�w��_i����Q��Lz~<���J�=ҵP��'�����/_H� �]�7Tj���2V�S��L���s��a|Y�ֳ���VhL�uZ�B}���s����&{�#�^��D��`�5E��\����Tsyx�M�.I�|1�s��G�*R�ȸ�bWlm��������&�j�z���44\ש
�q���,@����ј���VsW3��V�ޭ&W/�X?5��0���,%&��(���w�h���)�M}S��|���;0�C룚��p���ٰ�����{����K�+�z6.g_	�HJ�N��)sL�0��~�8������=�O��i�,�?���988趷n���AxD���|����j�������ǎsչ�|�)$��B}{Y�dK����6'|�a��(��b���	j'�a�;U���ջL'z��M�yRP�+�l��Q���$�S��lu�vP��r?�G��#v(�},ܡ5�9��O�U��MA�
#Jg�b7��Q~I�`���IHe�TS^>�Į.����ܽ�c8����nc�@<��L��ڇ])�Yx֟ߴ��V�W�\s�+J�:b��vq`�d-���
�_{��rt,pK��jqq147Rq3k�ZS��$cAN|#���~�|C���#f��n��/����SE������VHI����/�2X�菝%{t�Z��L�1c���4�_��vF��i\�s�����E��Y�͐����
���\xډh/�$K�U���iERu���S�9�o�J����vNjy}Е���\��ܐ�"h��$�yuQ&����6�1w�j|���>�i���2L��7t����^2��5X��i�k���<]��E<��$^�,���Dj��o�d��?�Xt�����%������[�$�t�X^^�]�����:�{P���(�N��>��#j#��I����V��G�½��e�Bd3 N�=΋8�p�j��z��Q��iaa�;�ș�L��}?���4��T֯s��t'�A.�k��������҇��p�=D&'2�����Ya(��S��b=������F�7���o�KF�M {{^�	��)����y�t��g���{Wk�>.��@,<�l��Z �4��f�*X�&�P�9������4�C��z��\}�wNT�S��<L9N���
����ӡ�I��y�Ax��újb���.�E��J�}q��e3fek<+�{-#:��H{yq@����Vyћ���KK�A���`�6��',��� o��G�KXGlw\Y��4�7���yw����% ̎ﰀ���|MJ�}����\�H�؟Y����l���I��a�栺c��J¯^��g�|���h���L��p,�S�v{���q�ē7hA��
<lm�R�H��wa}�c�l�b��VAn^��+�}��Տ�qk�;��V��X�
`D����:���������BrVS#��;B�L�i�  �9(�:��Gl1����T������;(h�f�����	I
�u�����}�m�~~=؃t�:O��i��&��&�bkq�D����hԪ�˟�.�%�����8֪W�s��A��+T�K᥅�[���FY ��w�F�k቎C�o�IL��U ~"��S�D��wu����T�ء�^��1W@��#3�]$9�T��s�1F䇸���m���.��F���.\w��P�������1`�L��t��'��"k*m���pY�ć8�����U��0��6��=�;�]]]���$3��i)�����y�8��=vdh�q	��xI�cG�&/E�E@^������t���0;�r_1Ҧ�	�Q���ϟ/ǲ�&IL��oM�{
��L��u�7���:�+�[(���ZE��DE�W4�(��'�5�{w��}����`���:�A�`M�΢��>@U�W�G7��"�3�0|\�e	Px���gk6��5���`I+�2�~Ocg�M1+����EW���E �����ee��4���,�c�AAA��j�ƈ{��i�$O����|(�y�n�bbZz��B��Yk���{�e�w�������<ǓJK^�VK&�`�1�S�|{�Y2�Y�(�c��mV��4@p<?�֖�B�F%����cv_�!�iLP����W���$ɂ-|gML���J8T/N],�M�d7�975t��|W�<AqP�d�����,f{�n�Ch�=�W�_	�[#�^�����x��ڀ�;K&�І��胣mj�!qw����'~�dwc�7z�A��ބ��t?��	�M����@��T���y�M�����FZ����i,�����(�p �����
�`�C��'�_|(X-���uh,��Z'�?�ځ�L~t�W��o����P���)�qO��I+�(�ơ���֥�ܒ���~�����lУ�����V��+�ż�8����	2q�)�Ѣt.eQ��#gqq�y��Kz�Y�= �P�6�-��5�x��OPk�����R�>�?�X �ޚ3����*�I��h\ N��Y�������ej,UY��Ej̆�aް�?tZn��k�^����{~�Z�$�P	�'���}�f15`�j�ܯ6�!wI�,L����&ͭE@H��=B�g��3�w���[�ߏ\���I��M6
����{�H�}ë,��r
	�:�m����% �Vi�\��1m� 饤���"��1�r ��y��Y��QFzlll�VD1M��\?zT�K�������H���)���iʈ�(;h `�Pҋ���
ƹywd$Q����mO̗N�z�y�u��2�V�x��?�\��m�����װ�s��Idq��;�X�֩8+>0�u��uը��Y1����p�U���-��
�C�8��j*�j�<#��V.���_���A��i����p��~��LC��6 0O}Y��z�}*/	s�4���;�q��I�wj,�4�g7��#I[��~�4�p�c2U�������g:7hH���c��<��׭5J�:��܎�}�}k�B4�Z��N��CXX�=�8�0w=1��P:MP���Ly$Ǖ�_H�v�at��g3�|3B3}� 3nu�v����ş�n���c�����z�e�6|�E���:��q�i�������I�=�ܳ�M�?L�ݥ�4�nB����������ا�O�_4�M#כ_?���tni�I����LȄ^Y�����3s�	$�;�����̮���m9c�^}�+�����!��̏%!�`����c�@��iٷD_�k^c&l�������P�i����*`2{���!%Em���Ƿ�K��S��UO�?��^�";�����H��AB�ev� "Cw:���\���q��<�_hq���C<9o�oU�0�W/Mq���>�HϏ����B�8Xǲ๗���cθ��2���߷�Ӑ�8 ����;�.\�RVQ(r��y��-HpW#U=8�N��a�W͛�Rw,�_��NM��`��@.�����<�SK����7a���BW�l3bM]P� ��ʇ����H*�9:+��j�nma�������ќ#9�a#e���V!�HVh ��l�)��I�u�<3�h�欞��Z"�rGxz���zM��}��e�w��Ɏj��qq[����D�C�2�� CuO�Yw��=�;}�T�R��fT'M�7r0�ڍ"p��^+�O����܊�� ��ݐ1>�z=R �?�K�����(9��������~�=�� ���Z��Z58|)1ދ=�:֝�N3�y��D9B�h���K�6t��ebT�?Mw,�l��JH?ށJV�q�^g_¾
_�QW%ïW9A_�=��9���Gr��⏜ZB�q���9�)�t�q�F���:�z��]d�� _f<���xd�L���>9��a�Dg�u����9��CVV���
v���i��X���SfC��U��a�q��Q��vp'q{�\�%����`�Զkm�`�����V������,bGY+?�-Z)3�3�^�(�
To}�W���No�x-=�x! ����|P̓ӄ�H̍n����;�`����:R��9��=e՗�o��q2�܅��𧱛e�	:J{���+�Q�z�i�)G���!���Tx���v8h$;����_�ulz#m���`|v�M�B�v�d�_��w��f3�P>ii[�1�M��'���.<R,�����;8���H%�v��<���Je&��1;��Q0r@��eH��T�sZ�-0��s
��v�r�fOʾ'��C#�ʭ�Gj�$�(s@u�~KZi.��e܅�^!�f�,�W)fV�c�V���:\�a�	A�+j��G}/0��m���x���u�,���`��J�4����c�������=m���
سV�S����=�\N(M~Rom�4Ec{h �`��x��"�6�Ǥ��	v����z0O�Ȇ>xꑦ`�
wb����]�A�w"�}q���[����f:�O�o/��3>�;'G�<�ä��z�T��5��h��L���I���e�e��>�����}�����di����2�w~��/ѰA6��~�����]�!S� �������&�q��ٓ��	B5�_[[�c��N�DPa�)Mǳ�v�Q&���D�_Fp��i��$SRR)��b�yz4�J��J�(��@�f�*C���D��6w�;\{{�Q�zV���(pG!x�d��E��o�4m����>�}B�1�=<16�.�Df���#&���vRVd��h?��b{��Q*��n����C����¡��������[��N˝a�h�T6��/"5���5
�geE
������ж���~~���&*J��~W+�Ϳ��$��KѰJ�l�����9��$��ZwBr��<�����HZ�s0�G$ �p9��#"�?��� ���&+��Hl�c��G��b
±��b��Ɛ������� k�4t�����Sw�i|G�um�W-15�S��G��Bܜ
Ǵ���	�j�X���,�r��j���� �*�@���jCi���n@uo�v��"���~\	�ng߶���B�ڈs-`U��oa�18?9�܏9�W���̱�;� o����[���n�B�nV]MM����^��l�����klJ��i���3�h7��n��3��Ʒ"#��r�2еUw���z��Sl���}�'�(�<�d�j��3�{NV�p�hhdȳx=���>��zr�R������VHM&`ݣ�N�Ed�?� ��&ѥf��2,7���]U������b��	���T�%�]̷_ɕ�;�?-C6�f����u��WV�9���؜�1�{7Xk�*>,�~Q���$aq�j�\�Z���:��s��)�����X~ԯD)�k�	�-V �r�T{�4t��C��%H@X8�M������"~Qz�'C�����S�I��e��|�=�_��޶NCy�FA�b�r˗>O�e��,z�D?Eף��'L�6��C����ق��$OҐ�!V���m.��@w�G�~���B�C\��C�#,�@�LPZ����0�v�T���R�P�PճR숵�raf���{�5�e�m�u���,��`x�]�P�A�i��E5��4,ߟ	(Wq�J/=��~4m]�U.J�1�+���g.�.���**M0Z�u>�s�$՜{���v��Q|�S#��پ$L�V��"��*�q��4�c^(��~' �N��#��8�*`
���<6�|���p��n�+��7`v�>4���0����Ό��d2��lÜ1�y3{��Wc ���O����JG7��/���ן֝�BbG��a-/ŝ>��gl8��'u�N	4����~��YGYA���WQ	���H�����'��?�C�9���M�ָ+����r�,Y�n��'s�,c���;���Ii����P�R��������$/��N�>��Þ��h��b�\Jܸ>�l�?S���(hl{U�qR:$���ׄ�����/ߟ��]~.�o�u�Y��"�#m4��ۿ�JJ[�nG�;���^�HC��u��~E���?�?2��,G�$i��bnͳ²31���s1]��<��hV'Ʃٴ�1�l͙bH�;j��t���B�m�_���Z�q�O��1�����;׌9!I���Z�"%4��M�Q���m.K��>?UvJkm����9�#v�agc��[�IWCC�k[�޳z���[>���1#��xƥ�Z�2w��J�kb�Vv;����.��rxD�l��`��ዚ1�\�3OA�ZZZ���<�I�=�Ex6;%� ��娞�h�8[��+��%�
�����;s;��|n>Y�� *�VMu֚��p��8ދ_�I�7�!{ qw0���SڥN_s�I��;�����阎��w��i��g.*"ۮ����]ŏ��Ȭ,Y˺�]rv�AlU��������w	�o�d��׉*:��bM��ݡ��k<�A��U���e�j,�z�t�3M&�����Z���ߋT�N�ɲ�b��W$�RW�%?��ԼH@���|�A�Gh���py���������D
��]"˫�ulZr+���H�s�T��1�ϥ8OrM�7��%�'�5:���^�R�!�@�����{f��2�����£b��Q�2�ؙ$ҽx���g��)^�ڷ�oy-���+����Í��}�ظ��2����$9yx�cBk�p<=����m2�zp��Q4�
��}�ݲ}�Mv��o��$��;H�޺����i�W��S�����T��_���ꣁĝ���`yi�f��cONs�����Q��snL/����ͫǟ<�Os� r i���훂�������4j�e;�U���tл���ɋ�#h.�Nc���:��"�axdda]��:���n���4�uZ�V��8�"o���$4�䓡���r��KI�x��_|�{��8�aw͔S�%u����S@��@yh��a�}�?��܆�z�F������;g�8�;�b�5�� ��psn<���Yr4;�U
ܑ���g{��Wq�֨�����)_|Gl9j�FǷ�K�+�]~�|[�L��p�ߴ��ڲ(�������}��.���ut؟z�!�I��-A�	�9ո\�碣]���Y[snyYJ�<����W�a;�*��\�@/��Ų$����yO��@�O��hh��Ԍ.�<x�=���@����I�Ʌ�P��4�i����/�?�; �of/�~����³���xGkg<<#b���caa![�bE�˫�vw�hM�Լ�s���ҡ����-���R�q�C��1�3k2��@,��� ڪ�2s�=L�5�\������s��(�D�	��n��W��]��n�r#E�M}���7��ݢgԌ��:��
E)�����ɦ@���j�������Uꂀ�*,q����2S|�>y1,��Z��S�F�S"�c�4?t�\(����s�%|�S���o��e�9{Ѽ� �^�y���˧��n$(/m.�As�S}Hb~�}iq�,u��������V6Z��ܳ�k�xf�mK��aWeh�����wu�wR�If��P�Y�Y����0h\����Qw�$*���)ҰA�]c�0��%��"#��F�k�8?8%�����3�����d=����j$ԔʥRO_?A\Bb`` �Er������f&_)�L!�=��hydYHn���~�M����L�ؠ,�H%����t`�?Xb�Uu��� �ao���*��;`K�!҅�g�2��'s�sVK�r�dC[�!���V� ں�V�Z�K�H]VV����2n�K�ݵi�H|G���4[�ᶻ���oc#���>52�51GOE�kfh���2G����޿�l^u�6�ר�����I���Z��ighJ輻�5�M�;���:�Ö�g�C�vt���GJ�l�� NN�(�<��+Iv;[oΏT`������ʢ�Q5����؞d�[-9.6�\�Q���Zφ�<��������}A�����=�B?R
V]��5 � � ._U��fݧ?v�)�뀫�bԝ�216�y��A�5��ţU*$n�gn�`�����իW��� �L�R]s������4��S������^�e�z��PC���?��x��Ĭ�W�����@֧t��d��������!]	7ln�`>{vhE&r����\�c��'��8�"���xp����&$FF���K��=Е���lii�T�*��H1z��D"ָ��F�:�QW����iȹ��GETz$�X.t�l�Տ�;>�g��+��{[�m��2��A�ZZ1}G@�e���YL�p\�* �H����׿U�1��\�^���*��׏*ZV+k��/^�---}�"`���kL�4[:M��QƝ7}�����َx5����<'R���r$'���Gs����L���Օ���L�S�!S���v�_�C����ٽ���k��me����6NN�GGGׯ����y{{;���;���$��±�[�� ��a#���J��o�Xo@��Wz��**7�o��~*(,tݏL阅���>5�,f��#!���߱(��\6�"��J�3נ֦�;�X���Q.������hGG'''�S|�#"�/��P�-��h����j�c�S#��6'I��"���Յ��KE�Y��E�#]���3ϻ\u蛡� ��F���G�����������9����@��N{�Lm#���5O�_M���ڊ���o�z+��y|�<e���G,,����n\��zf������T{�6��� �o�����j��*oP�f��N�3��LÚlG'p=11���1�=��W�͙�4�a��Q.���_����P0z�{O�'f\_����
��:���\aG��K�+V6�8/�����;/}��S��N�ٙ��?X{�e���,t�g�{��"�M3 +�TT3w�S�B��-K4�@��Tn���o.�Z��	 Y]��,�I�טE\�������w�xoWd�5���s���㯞�����7Z��"�>��jGˠ~�u0Ah�k�<|�^.T}&�99O���틞���bb+c����G7�O�%^I������@A?
�/����L���7�$Q�GhM�Bگ9F�]��PhVͻ}��i
���m���1;~�������6�c����:N�=�Ј��� *
J�����}o�EU���JǉTp&��ǘ�0X#<)�}�d D:�x~��u��	 ������T[ϼ������6�BXR�;N�${�ul5�2����<���Y5Z�����Lb߉%�9ɩ�I�n7k�j����sI�+����'}�BDi�q����� �z���aRBZJD�D@Z��F)�Mw���l����DE@$6!nR�- �����|��k�sTp3�ֽ�{�̚ƽΩ6���
Q���v������Y`4������`�}h8�vw˵���y�b�����!�A��d�d�IQΝ�w�W��<�QG�rEp-ź�eIA�w�����Q���%��-����E��v2��;)��@h����/��%jY6Z�X�SW����Z��#GI���	��k��Q�v�9j��z���w�T?�W���qE٧�W�VW�n�@�F��<�)�(EI.b�S��f�A���k%[�"T����u��	������C�\�5�P��,!
�$����ö�|&���R�>��m�E�+�&S�ʕ��ҷۘ�	�2�<�dx��gp�R��oVW_�a(�a�䗾>6^��y��D!|�!�]��iC�'��f�5U
�6X��좏����Rj�q3s�����;Wάx�%Oj�2x�S�M6��������K1ҟ�73�j� �[�'�����tM�"*TZv�K� �m 8���\R����5j�(r���A.��MjР�eM_w�v�*y�p�\��"c���M�5�����g��+,++S�=�O�S�1��T��d��]Ac9Ӏ)d99�_>݋ �d��$�0GX|J�%��f�kuI�R���s��op�ۼ�6�֝�1��Kb��갦553����˪�U+���ګ];��hZA�����^(K ��r���E���2����X�^k�}��WcQ;�)w=�P�:��J�!�u�3�fNR��.�vnߍ��}Ĩ��#^��=����Էc.�!��X���)�و�n����u��+vŬ�hڝ�R3$��G��Yӥ��6�����Ư�����g��v��8͊��Zo?�a��*D
�B�+�*T�z�EĲc;�R^n?U�`͔�h��@�kG�$q�ɓ��N ��K�@��Y��<��@��ڐ��-�I�a�r����s�s"��[�a��Z���;�T����+���gR˭,F9�w��x�~r˃Y�t�pB���l����~�:��p��/K���*�=G�vM���D�][L���r@tf��y��%I1R����`!�7���֗0o������T J�{v� dle '��kl\.O�k�E5[�t ��ۨ�ˉ��z��>(�>���ш�����������&�TT���*��Z[���d5??�$��t�p!��epӊ:�/�ֱCb���[���[ќ������r����Yf��g�~'��ss��*O  -�0�:+�<��Z��^�oOOr|���z��;0%�m�����|��T���ד�/���d`�`�|gyhUQ��AHD�
����{_X��<����|��M�i��Hz1@0'���I��~���-6����0(�:����ݲf�1��'`�x_�3�%#��D 3%����ˬaي�~�i���F@m%ɎC�;R���p^�Z�!@{g�)Lbq��)�J����c�R "�s�V��C��0Ϫ�m	b�/�@�@�@�Y��n@P5�.��cT� l'�>�4�k��'�W]�v�(���C�uT�j���h�ܱ���ぐ���S�����!�:W��������Ӡۻ�V	;��I?;����5��~q�J��"S��~󴰑�A����P�~E�����o4P| ��=��m�N�ΐ�q��=8�V�S��k��ؿ�зl���v*�j5n�#T�ǩBW��Řg�Vpp`m{���k�'��ME�}��.�|��|�w؍Ilu�s�䭏x�#o���:�]�_��'l,�
�M#cɺ�+mv��+2&FA�0���v�jh�@�14�]������U��"�ⅆ�0�q�<�oS����|��cg��B����	D���w�/�aW��������
�#��-�aZ��45����O88y?��8wnj@�q�؛�" �{V�{^�N���n�~�`�<���^N]kkk��N!���x����}��R��<<t�g�����jqlJJr���о�Z�x+2���n���eIq�
D�� E�c�3NM��fWW��;v|l� �Kߦ����u�(�nX˖�o���CJ�R�XY�2�N�o<|����Ttё 3�����@3��� �c�UH��|�MI�#Tc�-�f��#w������1�NV������I����s�Ͷ�U��ᇏ��Yy7(�M̩?��a�*�3�I��O~S-dz˨���J�)WK����
T��}�"�����A��s9jק��4�vIC@�ʁ�SZ\���L׮Q��H��j́����+4��g~˼�\�m�1�Vju50c���93��EP)'o''7>���J�2@Aن�[� JE��~�s�����ݫA�8�o9>:��=]�o�+��l?]��10� ��* P'�ù�Ӑ�W��ȍd���k�8~��P��Ic�����r��G���}[Z�b/��P
�� 9��;9i~^�N�Z�Ĉ��������>Hao����	��ۃ�Ji��Y2	=XW�wþV��q�L|)kS�L~�����9M���pWS�܃:���.��+� ��n��$�8���$�5�`������څ����Jok�
���'8g�w:T�?�Π˝�%j���4���N���F%�:a���ܬ���[^�n8|0O//��(����:(��5N2���3@h�H�;�*����:���a[��s0��Q�GÄ%OφF��g�J����? ����kV��K,��Y � l��	,�o���a816ZqѴ����v���)t�*
ID�hX��j�S�AK݃r���b���n�A���1�+����7@�4����yH�<X{���z���0�g����'rr�P�H������P���vv��߂ ��?_�Fz}��ȻH(3�'�d dñ1m����x��*���Y@�Ђfn�s��ppk�� Q�5�s�����KK�lɴ��׋*U��28S��D��%A��#���~�f�?~���w� ށ������!A��=T�
0�
��8��۞_�/�<7%:��IgC���6�Ɋ�'�x�2^T=ym>��r<::z۴�b���g�e���貇h�j�P����g��KH� ��RU�x��q� ~Z����M�c�
cۜ�+�υp�Gt���6>1V�j}��.}�]=a�I����Uo+���P���qPa :��1+&�~~���PJz��]]ݹ�O3ϑ���箇V��:�����w�! �K>��m^�JVRb1��llo7Yt���6��#�2X;>2���N�|���v�3�Q�[ݴ��Ő��k������H�B=�5eF{cZ�7f~'�b���Vg�^��[��)�/�{��[�'�m7^�[
�JP��<�Df���4j�lt��Ҿ�N�jg��D=�5��>���?��8�bX
X��_����C��b}������ �$k9����l�� W�B��j|_��)~��Q�����Y�ÄG��o�]��-Sa{���&�}X!־��KÕ�vxv�1�3�ԭCo�Q�[Q����Q�L���֏&TM��eٹr#�)0�~�~S����TV��2t��
�h�n�SqB���\TTJ� ���-Jj՜��.����-�C�4�7��D����"K�(����ר7n���X��-�OІm�����@�\\�A�����ly���� M��p��yoooh#U��)�lm(@�
.���t�
���
C�(��2��RΘ��Es�0H:׳��R����03\�]��Ó?>T����: ����3#ğHB�����G����-�k��TkkZ.㣐�AK�W1� ������oCű�'�9;�>&p���:70Ѽ�ϵ��l�u�B7t��I����ڟGx��p�J�:��%x����7��d|�	@�;ЫЎ@�I�K���EfV���I��;a����k�*����. ��������&�(���.w����*� n�pvgk��4G���wS�n��Uᜉ���241Q11�=�
�a,t��p�������&��H�AT�SκIL�]b�c��O2�s.��������H�4�{p��w_�������=?1997��' ��i?�4W���o��Z�%�H��#�?`�jy�<��+P����JaL
��[��*���ӵ��S��Nש���3_�?z��a'��������Rr}����tvwM��mhh�Ʉkk�������yM�1.�L��ӆ.��w�D���R�؍�+�m����%���'P ��6<C�끉}W���з�"��@SS3:]�w͖V�F ����!�XP?��j*��9�΍�c~L>�����m޺�3��ʻ��Z�9�o���_&�-�6+)+O��'���744uudffg8%l@����Q��ķ�6:���WD�\��ep�����6��P�V��R�3T߭��X���y����:Z���a)����5fL���0����8�&�^%̂��
m�9$>��cs?R{�s��V��ON;�����)��@��zQ���)����iv�Pi�2���c���ITT�9��옘�����������c�������l|z?Խ�qYRH���= 2�m�x:1 V�o�PC��$h����u���Z�� E�d�_������񝝽׸��'^�m`�:i��u���h~�t�C�L�?���։?��i�-�~�+�(�~E�JY1��VO���t)��/m׷�&��P`�ꉵ�@��_.�F��r� �.}ئ��o�%�@��@�yk�N:�k��]y�C��������k��0dB|k�6e&��~7sM�����N9 �|9�q�2��ep�ˤl�����w��b?�5.�S�*@\���_�hR3�T�����[L7?������r�pw��D|�����S6?1Qt?pCy���M��|�I��X�f*p3��o���'���1����.p������]��	�'u�ܱ�����3�Y_o��Hl��c9�Ċ��|q�A:��Ί��]���c�{�`rS�P�SMr��ȋ��,ǋ�Ϡ�H�V�!�U �omm������p����:A/���d�y���Q�F6o��`*���ｑ�(�X���dn���������9�}Z�,P`Q��
�� �;��7F�������B<ζ��SRRn�(�������c��%;���ڀ��Vș��Y���6�p��oRp�>Z�@D/���a�kV�frV�;w8ZעWƠ���<f��y��cb�=6��W}Q�M?,8�h�HB�$u:6��3��_x�*���ԤT�6��9��A0���]*�`�T��h�����@�3�r�@�ж(\�f�̪]�!N�bv?�I4���5_���=����v�T�.-��s��1����9?T:
�Wl���5D��k�^Cc#�U���Ufqfff=��fM?�Rg���#�~��lvՎ��՟���t+/��:��G|�o�[���!b'k9}�=�eU=c��j��Jq�c�X������OLOg
552�1�����=$*���K�$���Q�K���)޴�՘/I��sT/:UNUxz$�?�377E�B7��VsTVX��l�jG�������g���sq����[[Em3�sB����:&��7���Q�9�C�@C�p�j9:>V�C����}��h�X`Qf��c����<��Q������ă���\'�4&���������x���ٽ�1��h6�w�ޔ��g~�����߳VU���7w
E\�5اlnn�O��h���@Y�C�Tyi�F<��}�ZY999�l�G���O"��%�+�F�摥cG���T��J~��YBozf<��Ϙ�y���3�qkL��烦��خ������2l��oSxW�f��������LYV����V�%C{���s��s-E{���A+햷�8��s���S�U��3��������+����%�
�''g�R���үb�%���:�f���W#��[NMƃi��z^�8�M�CM����S}��FyAΞ�9�@�|ms`9�ҿ�-8V�^t���Zƽ��Z�K�΀�9Ѐ]9�I���'}+�g֙ŀ���+�f��|_q���*ooG�Z	�..."��\�d��%�3�{�z\-���yҜIݰ��6��$��g�G]���iT� >�n��5����� �yG�I�߿�<�Q��q��z~

=����i�j����7����Zo 9��L��n�_�o?�ӥ
e�Q�?�z0I�G�/��������eGkk+�i�Q�ؒ�їC�[�}K{�4 ,��/�ЦU.H��^gr�{���c�����=�M�T9M�3�ͤf���t����M�7\��j�}5�����a�䰵�uYU�V��
=M�T^~b*�b�6z���/W�gA�y�;��`�'��4z���i��Fa�D����z����˹
��1C������,-����Jf�(��"- )7Vc�����[;�g�g����:�lub!ߣV$ظ�0�z�{��-��&�9'���ΒQ24J�yZt�>��12���;cE���2F�V� @n��Y=	�|($TVS�yu��ЕE�[��ϙ򦁥�:(S[[[�_H�ek[��@��\(&���[��@�Kl凜]wou��!��i�<��w��\vB6B�xn@'��HB����^������b���aV�Uz{�C(�\9���KU��
��+���u��j�|0+�.q/���B�k9�����:݉�!��ϼ��Fr���@���wa���u�a�m~vw���
:ϵc���F<{_P CAA��� �z�8�)h`J�uZ����p2@���u�+ukM[��<�6V���UX��=�J�?�<�)�M�ϟ��@�&����r|���Q�K>�-�i\�B.�"����$�=�	�^~��Dl���,^,�Ie���}��f�|�V\�	�c0��گi���ܦϋ��KoԸ�;�~�Gi^��~�|��Xс;�8 ���Q��� I�Ф9�^>֘���>h��P��ܝ�����F��U�p4��cL���Qٯ_�b�KU�7(����By�:�T2�s�p蛜�w�?����Er=�)3@oAiv�w��D�c@�{n����������x0j�eH�4@��ԋ�ܜYx��묟�ƫ�R�F=c��;D���r	��t6���j-;�q����oҢ����4ϣ�a��U�۹�cS�`Ri�ݗ���� �)|�R��~-W�n�5����(��峺�v���s�%k�"#cc��k\B�l��s.�l�c�8Y��u*�P��.~69�[�U�~S����9�V�d)iiPf ��;*��l�A�//%��-�	��ß���T6�A5K%v���6P����A���ZU焻R.���`�w��^��1��!%�c:9��C�	���CE�T\��rA��ކ�5%�Q2�������vߣ8�?X�`t��*��~���dT|��s���
�CpnJ�bod����z�D���4��$BMB�
�O��S�UM��ߺ��Dn��p�z���籢~pj���K^�NqT��z�	)ݲ�����.z�Ey�辜4˕�k�x�5a����5zU1�$�=<t������XR�L ����̲6ϊ����蟼?G&�WK@IFūA���b�&��F��*��\�m~��~��xQ��-w�o ����ٿ��V���v}Lļ~�w��v;kț����o�:Ď��e�5��@B�7"Q/�h�J3�["�Y��M.��_L�ݮ*u��@6{hp��Td��_�D�Ȕ�ۇ=�������⟘ӟ�*�\"l���J4��a>�ք��mU��G[HaM�j	*�ѽ��_�����34�̪�ǰY��Vm]gb�tk�6� 5��?�_�]�'��^���d-����T���L1wO��Re�.�T�p�K��Wm�;���~��GNp�f2I�����v�t����ᗁ�v���~u������ÒH�ƃ'DE�ָ�%�P]�j��0L�1��~��D7�J�4�y}^rU�wf�}跲�c������˷���z1��\Ͱ=��	�A���BϫV�]F���e�}��m2���-���kcb�V�%���0��3�(�m�4������i��#yM�Pz�������԰0����kվ�*=�j�P���sv98�#�<��O)mW�w]v�G��5��=�\�7�%����<;ޙ�@�4x���C�c��� ڵJ�{KC3����38�B5�rļ9�v�Mf���I�f@Z��k����*��8*��d������1��r*5��0tJ"pbzU�8##��㳛�ț}|��e�w>���@y�?]��/J��Vx~������[[�|�〭A�^��`-/�l�}?�>�@����4��J�߉a�7�#W�ԃ� d�*�V���P�by�~ˈ��~��[%����ܐ�7�z�aA;݌�Ig�W��j��6�ʰ�Ȍf���Ub�gvB)��,]��-h{{n^�!m�ʔ���6����������+��&�K��m��J���K���3��_� �֐���qj�l��9�߈�J��S�����Br��V\����@����i�o	R�����1�{h@�C���������V���gn�E��ۋ�r��_�SǾҸ8���,\�A�}a�W�ȴ����u$йPa49��;�w�)P[�j�4V�;��=�vC�83�d�X$�t��4�m� ���''�

*���JUq�����7�;�����E���n(��n+&I�#0۩~�����>G?�VH�qO����>�
1�?�ׁ�K�R�iv<|"��4�ka"�8��z1&6Q�(EI� K\h(�
�O�GԒ�V�t���K�wrw��z�TIݶ7�ᨋJ��O��Nl�yLOm���w@�x|b��r p�&Wb��4A��0���q�ʕ6�2X�����t���@jL@Hkjj����V3����ѱ�O&�.�(�Ǯ"f��t%"�ľӊZ	�?'�b=�3����+�3G!ۼ�ڭ�Ɏ�S�c���1m�Pxm��cgg�5Lw}%~
���}f��Ѧ�;����iU[�Y���v����?A`p����C��;8L��U0��ƮC�rzz魭-xU�_��}9�o� ����2u �B���h�k�x�����`�D�//�5G�{���bR�XG�)��i��p�f� ��F�����*w2_��ZUg�8�Z��� owv�~]s�����G�EZP
�����&D_	���϶^��R�;���?A��7�|_��Q��<����Q���W�cp˻}��w�Ӛ���@R\#������ ��C��(��zc�||v�z��C��R���7�T��z�1_C��^����7wϯe��3N���[��w5Zι��Ҋ�A6���(��<����{�H
�&�7��:��O�/XR��� ���ŋ��A��&Y��?�҂<�7ea�>jr�i.�� T.b���O��q���y���4#$$,���pa� ������<)��ќ�o�m˞�6d�ui����R�xM�~�@+���%��"���t�>�V�/�lŗ���Lڶ���n���]�R�y�g;kj;n:�E�c�Ꮵ;O�Sé*��ٕ�|��k��t2n�sH��Y�W�tݔCf����.ccTž8�#%
���u����x�k�μ���Ey�O�_w��կ�Pl��;J"x���[(��6ǳ���?�r7���'g����ߘ��m�93���L�-;�؆�ӧOߨ�zušZ���)_��bzܝ�r("	c�-�#�W���sg{��^9�Zv��-RRRBF5��XkC#�����j9�����F�P*1[*���bS_��0�ޠ@�m����L��fr ljjj��g��uj��&�������c��lpn������_Q܃g��Ni�d�T���j}֓sC� ������k��S=O{��"O��P�msZ-�H;��n�1o�)o�I�53^ll,C�
#9>���e&�RY�gƲ��{7%ɲ�PK:��t�J)���uT+�h�OM���AC��U�~��m�������kW��֖_@ ��/��#�O�/E�\E���:&H(��\��>I,��UQ���Y��Ls(�=��J�R�������i�\�M�Y�~��e���A��~�t�6�!%�L鎂��vz��g�m�u��mCرv��T�`��2m��`�5۾�+��1P0�1��� ~O�f�C�+�*�H����V�n5+"�a�e��F�+z��]�ӹ0�X�Q˾�@`wA��n�Tc�͉�!��-�ҕz� aI�\O�������Q��ks�\$�T����b�<=��ʺ���~r�/Mŝ�bV̉��n�ڢ�ĳ��Ӷ�y�ć���?-�Ҿ���W�.p'|�{�;xCt"�$L��r�<ԋ�~��\��N�~��hy]�g��A}���o�����a�s�3�n%2b4x���7Zg�665�ttZ���O�#}���(���/��R�f�!h�~t[^g=B��d�'��_ؾ�L*�}>Y����0~�┑9���X�YE*�KO���-�_��UFK���������pS�"����204�98��Y1i��q�vh��Ko2%�<��=�An=�� 1�˖�i��f���0l"C��]F��:�g���9�К�>{�7�$~�	cA!i�e�<iT�i0�p�!�I�pO�Q��x%�'�2k���զ��$�R�YxVz�����
BV2O^��PS��Y4Mp�T��7�q�{�,�od��fTIiT9�$�-م�A�v�mUeˋ,��^��`ꏞ�����.{�`NF%������y���z��o�1]��#��"����9IhB�»S�S
�I>�%�u��A+���9��f���2O^��˻ h0��V�nX<�D���o�
�Ka^�ċ1����>I�{WX)�ݬ=�]���^z��O�w��}���q��!o�fƵ���b�"�τ!��ymy�-���� >�*�W�X9r��e�����\E�i�\-)�_|����>������=�5����ig2�z/���:�1��+O~la57E{�JT�]�sX�/ ������:�>W�vW����Mے��
�`V�<'.��������Kw�����m��&��xF��2��J�zJ���]N���N-@��0�����|?���#ؗ.ELp��;O5e5�[�Z.���".:�I�
��:<=�{G��:��p7#��`>[צ�X�_h<��˲k;��RG�x&.pA�]�U䎽�Ӫ�������c_'����M뼊dV�s(ܼ���(��f�a�>�Jmd�Ã�!}��m&�t�	�ӷO���e��'�uu'���,��������f�b�_T]'�A���@��l���I]N��x�y�'���
gN�u�����wI[^^�o杻���ΐ��v�>��j�VY㘭���=��c�Yu��nAU��C��.Ů-��[�n���K3��Z���0d���E���M�>�/��T�ݐ+�#���DKg=)��ʱ���00���ĥ!��km��8�m��=�B���^h��=�}������)�ﺦ��e>��M�T�4��x�H�_X���#�=1|����?yZ���H˂9ʲ��.*b���z�H[[[��
��0A����0Ѹ���>�ّFˢM�u�n�F6�����w
��,F� q�ɻӁ�C~���13c�,b[!{�|
���~�]���Җ������)ACG�zZ������o���b�Aھ�uӲ��҅��=QQ�M\���G2_�hlo#7|%v�]Ò'�{f���Zt�I��L�����p/DW�V��E٠���ǟi,[`�;��<�i�#ɚÝtg�����i��b�O'��6C�����Vr�ӣj�-�H����R��Y[c� ��:������J���������Ғ܏�_S�Y/ϖn����V�)fWZkpg�������ݶŶ���  ����<q	}_s����
�tɨV���)J�'��|�{�9Ue�(	.���8G�d �)f�?��� هl�v����{r�`�Y쮖K�x!��H���Q<p����%���ka��)������;-��C��M�^t�|�� ��G3��aJ�&��b��H��j����p���3nv�7���$��г}�l�5or(��6��_`X"�B=ww�ellL}�v��23���Y����c��O+�i�@z^�}�ЫĿE����-ڀ?=8/i��nɼ5�tww�g�.�$t���cCKC�� P�"�R�9�Q�G[��I�^�z�Sqzyq�H�ENqߔ��(�Θ�Z�V*����(�\�ş$U��-!k�����ڑ�d����7�.*����X)��+�4̜�j/Q�
� ��ҏ�Ҳ$?�ׇ�0;5��M�ԛ�`��'���V�R�-љGeT�+[p{BlU}Rчe��m��n|�H^��J��O}S^�(��O�\vZ�����I��r#�֣p��i�6��ٿ�C��?qJ7)�{X���y��}�����*�=˕��n�w��H�84ivA��x_�d�=�rH�g�4���j�!4iqþ|�/$$t4��Ԧw�I�݂w�6��D=N�Wf�?9q�����x�/��5��2~ϓ"VE��󇎎j&Z���������j
�6ۻ���.q.LFd�2a��Z|���_��
p,�Q�Rt{�Z��w���{r<cn̸~&gܼ�[�Ўݏ���S۶w��%?z�	J��[_�q�_��d�h[c\T�y�q�`a�T���)
��!�x81e����B�|>��an��#�-�#�z���pU�ez=Fا_�m�ުZCwAw���r|�Iد yȑ6[I|��c�>ߎ��}G���n�3j��zOOE�J�Y���J�U=/�4���A��|�b����>%=n�������RVVnv[��2����d�.Ցʒk1Y�R���3�#��(�^z	1x���,a�J��x7v@v���$�.�2��}��M ؅��
EZ@sI�O�1nZ{o'�ƿZu�n�E��@B/��mX4�E���X���c���ؤ�� yY΀#i�,'����4��|�$�Ik��1b2BsW�HR�
4�5��Y��a����٦�5�"	�}/�H>fA?�H^�\��l;tz���?�6�u8�������p�gMz̚ԣ|�#��v�-���{b������������~p4��yUj�{�^��x��;9;���9�
�H3����ē������Y ���O��>y��	:R�����tz��YͰR5��K__�
k�ͨ��E���~�V�]�	ь_p���,�LT�@�t�m�B�*n�I��0���-Mw�88��q���Q�V���Q�^7���<��Jw��v�������P�?}ɋ�in�e� Ģ�"�05�U+�۟�����=�� �FC[h�MMM�P_�%��=�H�t�P����`t=6km#y9�@��o
צf��T4�KWQ]��ӐU-� ����b%j��B¹��[�Ehq�bTX1���� t���sIO�kҝ�.��� Q�OJ*|�	/N��v��M#���bE@P��j���i�Ċ��{�z��M-6J���Ñ�8���F+3���i9�ݺBL���������M%�o��%`��wc�}6:n�����e�Fm�`G��0�e��ý=�_�>%����Ҟy�R�~����$�Y���ݾ�5hn��m?���q<ck?[����������9
0�e���cwZ�p������X��1/]�>�$CL�8���w�4��K���3�ݕ����S���2�����#Tsgc;F�N�-MP*=�R���S�hr�ѫ?B���ho�5h���Y�1ߵ�ӥE�'Ѝ�h}�[?e���#�@K<�H��S�.����g��~�w�l�4H�[	Dd����ѝ�x�qy�JF	������4���w�f��o"��4��J��v-�5w|��mN� �� ������{Z8z�̽�a�������E����R� }��=�qooO���N܍��»��l��K	RDh r���Ax����-.jݩu��_�Z�fIF��w\�u�+9ő�4�wo��D�����T��]K����F�+־���4r$���T����L�f�z��~�bbܦ�] ����p���qC�ZbACMU3�(��Qc������F�%�i�i��~�◔�`���ˋ�0ͳ����Y������;��A{��kǙ�;˧��`����E)�jA�J���,wq�j�k��t7p�3��)RA���V���'E���6	�g;]	�KPa#�	������*+m��#R͝�F��U.HU�2a���F ��47�G߈ ���;y���Vm�woe�m��4ޏFS0"���~�ES�<¶jSS�k��Ѯ«��)������9(2���$��`i��}'_q���M����"wp���ʟ���hoTX�����|��J_������l[���~������ ��M�Շ��P�|���B�C?:�ٟ��V��/9eq>.�-���ͤ@F�+��wz�:�P�����9�y.�L�S�]>��0u/:�o���R��� �p&̞��.�r͕�a��l���u�)<ok�G�Q|��]ϙTzQ8�w�=_D�A����.c�呋�P����a��t��y�Yr�L�q��L���/_nX>����3���L�0ē��4��*K/��:55F�� ����m�Y3�.��&�;&D�|��������s��',ͱ�5!���j������������^]~c?�/j=Ԫ����^o0uR�Ļq��5?��J3�p���\���~Xo�l���M�R��Dl�GX��#��q�܉�g)��pzG

5
�jy�v��a�3
�5r$���i���vO���H��b�JF�e�>�����X��~��ٶ�}K��4��c�9���CԔ����wQ�)@#66� �<�MJJҘh�Im6G8>��Z�Am|{�*1��6+9ײ���F�^��ZMK�u 
����=�S����~�;	]�G���﯑��Aሔ.��*vr� ���@���<a��0�(����~>?w�k��'%�?*Xͪ>}��gAp��޷��#8n�h��z�$�/�5��������S��۲�L�#dI���.e�p{^Ua)���y��#��4;x���㛃>�]�m�?��@���*����O�11�7A��k٨�&���YZZ���ׯ�@����;���5w���5��VcdO���Nf=o�4������p��7�/��7�m��Ode��UF�(a�h�=�2a�~�<p[���r�|�*�������.�]O�t��Ԯ#�q��rȤ�0��0�Q��/O�ʋL䬣XP�/`|�J�g1�����90�7G;!P N�����#%N7�-�{P&_c�\��p�|β��1�e�Bg_K�k@*@S��k5k�bJT����"+�����-xp�rW0K�q�� �'E���Z����ڑ��S��࿋�3����A
0/�gN6
�s�~�ʇ� �T�+e��yX�=:���&���C{+9)a�&ME��A�p� ��@,�����#a�	~����^"�����0�b]��$5�t�I�q^�����ˑ_�4,�@��q&�{L�����1{yNp�"-���R,�4��^e�ؕ��("�u8pv��0E����ɗ@v�n���y��f?�$W��7x��-��(n6�z�ߴ�ϭ�܄!�[����l�C�ڒ��[^�Y��G<9�:g 3jk�cT��d%��X3�m��M]Pߺ/���d�����9b^���[QU���w��4��	��r�X|B؛�L�]*4A��.�)��W��=U+o#nǸ�?z�)��4�������S�p�ga�z� �ג�%�:Q~o �j���s �,�f�"D�4����p��S�a��dI�l���N���6�~4v��+i���l�ͱ�d;:��jB��0�P��h�6�D�ڌ�ӱ��z7Ě`#�y�j:;��c;���9EU/	-	K��k��91��9u� Q�0�q7@�	E��?&`�ilaD�%��2����[��H�)g�铙��Kǽ[��t)C�ϗ��S�c�d�����ƞ\aw��*����K�s�.����]�a�����	�	����9�u1=-��O �H��2v�_���F#S�	c�[��%T."#�2�v�{:߿��syq�;���9	�[EU���eo���,�����\X�I4��x_�K�Ձ���	�my�Y5B��XY��x�qw6?8�C8�=uF �����j���|_C���_a��D�S�Σ���E�7�r�|��rn�㜻�?a�g�)��E�]��2NAUw[����������3�WӦ���W�檛}�G�mr��7���p��2��mghy5E[	� 5%�!"��}��]�bͫ�.<�}S�5�����-���M:ڿ!�q14�&��
�"�S'UG�.��zwl�n��a�<$d!?#����Y����`z�5����E�����O�j������)���=|S�O{��v��Q������0��u\`�a���/1ȓ�F�y��J����O�rް:E���&�{*�bee���A��窷�B=����6��� ��-����0˥n�-�������Ĩ��KMF?8�C!��S�^�~�Ǒ	L�����둙5�l�l��(��[�M?3Og���[�l��~�wr/F?���D��\M�\,�i�<yZ�=�- �m]�{���p5L嗐:ޔ�ì��88ǘ�ࢧ�*1�%2$��夁S���kl%K:rjqZ�#=�[3`��_VD���ԡ7A|u�����#��Qү�o�]!?YO=��LH���R�7\�3���s��,I��ȕ	N����u���Fo'^��:'����miȎY�?�A�Hݜ
E:���/����q8y��K��.�iW�8C��5�������Wܼ������W��_�x�vǹ���.��ȟ
ʊ�7�F�/s�����\�A�_��V�/�8)c�c�%<��}��@s�S�_����?�aA�T��w��j�X�����9o��>���h3�r|O�Ry󟼳݅��j��x��KF�*�1���n�I,ݿC"�w�jM��KL��1k裠j�%A��| Ճpo���dbbz?a��{��d
'Mu�:�v=-����y�Up���Be���_ǡ��Q�X;gPԐq��9}�t���N1��qȣg@��#�� �E������Zn��=4L�G�z��9z�R;U/"��"=���	��(wFg� ��X�mX|_�6�{��B} #��y���������G�0�cX��p/���Oռ�iܩP�oݥT$����� X�!+�+����qj�4����������1���8�jÚ0�,_"�R���K������^�b�Y'u�6g���d�
+������p��}�Ju�� 'g��+}q����57w�9��(��)!�}/gE��,@�Wa�M��9�(�h����
����mA��PB��.IA:EJ��;	�Nii�.�����f����{ν߿��yD�k���;��c���n�P�V���j|�f�Q�3o��[��n�5Q��)���R��fM.|��=`H��nŘ�t"���4 ��*�|�G��Ls,�>�݋[�7��GQ���*��*�tO�Տ
����|D���K��9/��/�?�`;Ra�'.�P�ޗ�D���iJ�p}������c�_J���-��rw-���sn�T*��z|�[��}9cj����OP�ж繋�Uo�:�8�A��y�İP_)�,"	I]3��4d+�����nA�D�G��X�`tr�����_f��~ڔIs����BY(u�t,�%��Z��m*-�-)�Z~|~ך�H9������U��9�,E>��r8K)>�l��H��Gt�=�L(?!&)�����+P9Ej��,�����tZwF���^��B����A|��P�r��G�����Nd�n}��B�l%֒c߬�;鈙jqFҎ_FOA�E~��cR��x*�~�2b�nt��@�	�N��ӻ���k���X�
zlu�goh�V�A��I����{|e������Ajʾ�D�A�~D3���+M�E�3S����AO���m%�Zƹ����y�U$���ʋ���/7^�"��5 \�!:�*v�C� # �����;�*{V�;��%z�<�i����{�F��0&����E��'KQ"�����r'��1�'^����T���!"�6F����bxg��h�ɿ<Q�9��:�����J��%��X���̋�̋
ĩx���m|i\�G9�+9����ɪ�b�5߬�����OD@_��YJ�1�7��!�W?L�Nի:k	�g"�S�Ey,X7�֝�-�Z�g��;��1)+18��QP�q�^�+��j�\���w��P�O��5�����^��!m;�/,,��N�Y.#]:+'�<�g���I��7eQ�o���������,�0���R��l��`���Y*�F��e���󓮷��Ϲ�;o����p	m�u΍�8�#h�v&8)�����rB��Q��dkR��Sw�D�b������|�jM�Oj:!+�{F�����]��uv�f�_���ʨ��$�`S{d������#�v��X?LF�2�y^�z]�	(����ῂ�-NN$3�S]=}N%V���x� r�h��sN�4p3?h|��P��0恡����!�H�!��K���$�i
�ܝ��]����	�WfL��L�2]�9��=%�R�Z0>)#�R�S��䈼�{П��Bo]%u�Ͱ����8���wS�
��r���(���e$���p'�4oBV�/�X�6̼����{�>���`����6�3��M.���y_Jo�?-TB�1`F}����w�=~�|\q�9�&��B�B�HK�y����w��,>�Ǐ���irˏ{�}��[I���h�ŗ��~P�ex��"�]�����{|}�z]h��55E�o-Z�o�[����C�nP ʫ���Mȣ?iqpz��z��f���hJ�a*r}ٝ��@o���W����r�6m����9
+��)�$c+Ϡٟ�4�5�Va}Bq"��E$��Ե�&jf`�u�;���6ǌ#�SE��v��������l���]J�ٓ���hs^�]ى�Vz��Jd�N:�#�Z�GR�@�Z7�q�}K���������-U�bQz��$>���yK`\=�|w!��?��[/�(������E��S-��H����q���M�.�[Jl��yq�g�m^�xw��rr�l�B)�Q���鞢�ڬY���7?��H}c�U�.�n7ts�%�{з�[���J����b������i~��=�?�ٍ���'�"h�9�����m_�?o�񛴚�tR5�ҼY�i'Y�T��[-a�G�}�{�CN4�y�	��^���0���CAz�l�з[�q�����M�j�0�\䲋�-r1�܁3I�᧔�f�ժg����Ab����x�OH!8~��|�B���Rj]&\>w8ؠ�g��t��L��ֲ�6-����ѦxiQ��o��˺oM��Y#Qb7H�f��y����Ӕ~�k`���&��F�^6���:����#�C� ��- �\T��u��66e�Jq_���|�cT~g_0��}>L�e�*sX�m-4.k%�!����V�f7�l}���	f�ͨqy�����������R�g-�L���d_���˖���|R ��zw#� �y��Qv��]/߅�q�M*'�S����W�d���F�*��_�А.�ݘ��}aƻ6n;}H�����1∯A:@Aam�<́�&�{;tXd�%��s�����{�ƹa���9��X�4�cr�+��e�~�@Zc��ZL�鼝P����}q��;%*5��\:��'�4��*����J�����mٹ�� �t�i=t�_B��*����L����$�����O]q���! !�*$��{�qu�H��&B�sU���|�����V�1���*�l�I܏���_�����zC���S9x��I�����3`�Jy ��V�~ŜL\x���껵�sQF�>���
�P� ��["��i�H@�:@��� ���ok�M�[cߺ	F^(����5��Y�?��D�mlI_�joOw|dܭ��yY��A�[9�nC~�=��R�,��b�rcIf��##8999o4���n�^��o��~��-r3��B�|r;LZ�ݾ�8x[� #��1�#Q���t�*e�_�7��D��Vm9ݽY�'�C�g��+�wǟ�`W��0�o�NTy��s�7jp��`ﭷ��ك�򞅄�9]���b���f�����"[��y�f��ܭ�&{<�J�� ��Z�>�+3�,<!	���ߐL�<=͗?��� b����kk�%�ߩY�(�[���6(��^z��Ͽ<#�G����|�Ԝc�?�������Q���f�?{�6L���ð��
�G�D>��+�Lh�n��ў����֜�s���<�����������0�%>g��V��g�FFjot�`޿�����bB#ꓺ��1y��v1���)?�7x�yx�L�:���������#MM͟�~��L��"�jHd��]P���32Ύbb��>��Dj��֜A$�[j���>|��ya���]�
WW�.���O�s�|��i���QZ���L%�_���\'�*1�7*F�vu�͊:��o���`X�+]#>)�ml���s��X�ak�
��Uצ��T��_g��Fc8-_R����8ߘ3<Os���0�K��_�
6��4���]~+]�hh	oO=���9��G�}�A�n��d5$fܲ�����s��e~���I��-�a�^L��ubb�>�@�/����.$��پ1z����^�����0�!���'��\�x�n�h��x�u��O�ש~m�Zu��gл����&bA/�%�n���ޛn�u������x�� �K#�{W��~��9�� ��)j^��P��^fz�Q� �t`����b�d�$��]�����Ꝁ(��[cI=�>�>�`È���-�\�5�j�u�&�h�߫�y�.�R�������1��0�O~�?�vUa�ɢ�}�l����П|��5$�Y���ǩ���Z����a���l7�Wmyll�1��u���Ʉl&8
/J�B
��K�Z�N
���ОM1�C��8=�N���*�*e@1'66����L~����'����v�d��J��<�9�)�OR�F.�/$��&�2>CF��ZU��;���W�]GE1,��ג�����Vc@qJՍ�i�H��|*�����;ґ�F-6��27���$	�Z_<���r8o�=���L|����)|�O��F���f�ל9��Ny6[^^�ފ%�5)?�իW- ]c��ic�]u�^}�j��9�+�|�	~�E�_A��o�,)�M������'$�N�|9e���C
'�Ϙ:6�V���ԏ3�~Nj�z�Pj>2�'�����5�ϳk��WR�}3��++��J oD�;J���A�+�$�S����
ȗ�ΆJ��û��̓�>Zك[Q�)F�o�ghk{�fl�_�␑��A1��?��)�sl�� nˇD%��Rk��ʒ�͚=���%;�O�.7�D�\Z���A��Cg��q�Z�����̎;��^�_v���~5��n?�����tHuq�s-����2��bTxVkͯ�fه���5���4���ȷ��GR�(�+;�ʕ��(D��1J=��ǲ�g�U�9�.Pl���?$*/�ǆN�~Wk��fY�>��.:����^��F�_Ϭ��Y]�85� W���η�8 \I�,'�Ő#_��j��r��C��-�}����a�=����/F~��Sf�$�~/�y�����; %R��D�qӝ�k�����U��PO�Lb��p�{�wB�J��. v�φ����て�=흃�w���������J?g�н����Sa�a������ѿ,&#V�����0���f, '~}�`�8�)/�8 jV��.>���vz@:���[�{���㷭~�[ʑ
C��'@�P	�?�K?�~Hw}V��k�h�c��zy��u+����c��ϻ��U
TUhq����,��F��oo����$;|�����l����/ip�E��qh�Iݴ|�լP�����z��r����C>
"6iQ���g�q�>G{�w}��u���E����	ԣ1$4t��.ue�;P�!lU�� �F�t�<�u^�FݟU�ޕ~��\��YJϲ�M�_��;} �:d!�k�X�O���:�(
ɓ��A�<(Yf��x�/��Y���ͽ��_���P�����u쫻~\���	��͗GVל�����m-���n���A��������jam9��L�a瘐'���H���5+�{����8&ݎ��@��ϝ��K&��r����[��E��OŰ;�=\��X3���?v�M.��������0�~�հ+4y��Ed�f�'Q]o,-�߾s4 @���
�Yz�1a�� زR�-�XVV���;`�3o )�&�/�Է��㣥:�=ҧ�/O|�O�ؾ��Ea���b>������E��_��ϋ$<A�c���he�F�w�nB��98
�� cvW�%�'�������TH]�|[�\�g�.
:�r�����Df�+��8�<���Ӌ{mn�T�E�{�h��� ������<��x��)诖�ުW�M�� }(��q�?3Z��}|BpWp`����Se��fBwۘ�VU�K		��?��<	��SA�v0�N}���nZ��h���C/����[:�� &o�|�*y�o|���������v��k��_�&���P�w�P�}O�A��@?�,=��V�L��o��m���
-��ܽ��ݰ������`�N�ZX|��s!g{���Н����9%���_�KK�iAؕt%����n���tJ��9I�9%�h%����j� ,�+���f>��ф�����@��L� d��.+$��<3�4A>/�ߺ��m;���QY�FT�ڶn?�Ǘ�$����DD�?s�������KS��/�۽����Ĝ9��Ey���%���>C <,,,��#��O���8��'�ֿ�8��"���� �HuF���>�Ըu�Faq�c�r}�L�n��A�kk9�F�y+����T�ҩ��gAF�m�`C�$��Z�}�{�e{y� �X�`?�DUiSShQ�\����4ϳg�4xxx�/(��� ��o�߷��T���r�IZ7n�6Z�-E��Q_#�[m����]����t�M_όg2d�GV5�s���ǌ��4�+Փ�v_J������������洈�����:�N��d�� ���	߼���,!��ܶ���B��h9�Pp��ÿ�{�N�5�j�-�?m��\ku ��Ѩѳ�S��v6���fG��l?��M�ɻ��ܚ�U������ 
�dg��1���U�������-7���U�Tj�M�u�[���brb2�'l}��4���X�z0�����8�U�i*
�~n5e�L��NQQ
7��z��@�؂ss��7
뛛�e֩��J�'-�)��󥷶����o	�>ʮ
TN�9ٕ�v`�sKQI��n�<k���՗���oa�3��	yƅ��Yx��Pi�t����S�j�;m�#�Ù�����.�_���hj$�ߓ�����}��2>!Q4+���s)�#-����P}��OB����߀m���F�to�ȕ��)i<J�㩬�;���C�������/��mm����]����������qX��dd%K����?�����PTW'w�D��4?�V`��CS3��Ǆ����~U�|/<�c��������O�C����WQS3�np��G�k�4��"Џ�m�"3��~��
oߔl%���9(���f
N�:X�'�:ɼ�m�)#^�4y���G�%`�:9�AEE]��^�O�%l��IIIQ��4{ Z�{=��?<x'[DE���ӿ��$#*ټ�֯N����0P�]���c�����[Ӎ�/� {�ʃ��\t�grnd�r�p�y�U]�o�-0g��2F��R�ƠWg�ƿ�"<�~�ܜ�Jf2a�	U(�
ϡ�)�����PM�u�]xś2���DEQ�I��|��pܤ,���F]�x�]S��t`i�OI�x�����)�ŭi�&czP�����"y,wE����q2�є���#yʶ�Z��5��tt��ө��V9Q�׸O9��jsE��%�ћ����>o~?Ӆ�6������7_�iV�+��޾�N�R���.7p��Y9��~���� 	���ò�e����'�t��̀n�B@�~j!�4�V���@ �?%��Tڰ��%TǪ��c��PV��roB"��%�~�k�vQ�3���&�(���r�9�f�Ak��/G�N$��y={��|�w�;"�38������d�C�{ֲt��d�"�^2u-��55�D��n��L�K�s�ԁ[�����(=���[���hQ��F��ߤ� !qty�sN�+ǯ���|�<�R��ow��m-ҾB�A>�^�,۶�P�Ϯ��p�l���)tT����~���P�Mm���D!/O;v..��4�XFĚ�ģ��=����8Y8>UD���}��k.�+h^���e�9�Ɉ��]+�<i��:�%P�X3��F�"g�P������r*��6�2GX����fҤ%p<�����U�Mî����{���Q�ǋ�C�_I^���*�����!�V�i��h���kn����ds�d����,X�h���_���I��z�óU�`�\��X�9�mS� �����T;*�A����*2ى7J���ZT����@ l����/ϏW���ע%�N�`]�E��hh��Pě�������-Gd���^?�j��~v
>�6yN���Z�KRN�i7h�T����]tvvF/)Stx�W^�u�v��4���o���
u���F؟e;��{����B� WLMMm9w�.���J�̛�U44X,�?uHj�����o� �W�V��`vS�oh��Xt*Z����^�xdU���a�1;��ym�+Jy��T$ZK)��P�9`��[p�J=M�$�Ϻ�}>Ł����Y{����3=%��Ca�@y�������Z��,���MoOՏNM�T�j3�-��$!~�ў�j��hOF�d�c�<Y:��8h��p��6���m�&��B4��G�{��6t5��1:&��5���gN��w�c���k	d~u@��p��Ҷ~
Ec�]���.�99QQQ����f��!�U�/_f��d2�"[o�x p%����@��F�s*�L�#�'����4!�p�C�yu��m��e��$��n����wX�I��ן��vAi��,MEZ�C>b�Ps$38�(޳s���1̎����
��:�I��x>�b�Jy#�yϵG�h���b�P.H�u.���p�����T�[�⺍�j��Gͩ�KG���N��^��Ed�	���k�����Fv�%�Y���Ծ9 �LMT��o�6@ܤ�ك.��W,��0+v���Q~N���1��/�&F{]�o����p��&����G��s�	�'���:6�ݎ�<���ۡ��#�
PJ��$4:���A�p���z~Pf�)��c���f#��&��/��>)�`�=�|���)��r����u{��PY�j6V���1N�Bg����|��]���ڭ
�������I�z��ı�8�ס����D���ͼ˞�z��������^FO�I��pbB
Vt=��&���H�_ϋ���􈃟���̵`A�HSSS.	k����<���9I���==�	C�R�{���DYR�~��3����-���xH���Ϗ��@Hٝ��V��(-�N�O1�<�$.��&�sMM>3K���z��X����.f�+�b��N��<6�o�ҝ�Bw^@7�A�i�e�U�L�������{���+tbד�����S��4uX��C�A�\n�AUTW2̢||dr2�Œ���FL�N����w�J�c�<�",�����Q��o	��C~f��g�xA+�Z�3I�lb�Ka̰:5�1���8qC%X��絍���cR�ۄd�?)v�n,��,^��,i9���o"Oe4K�Y�a�QTEE0��6 ""RQV#�����Dz�g��$�|UUUt?�Opʀʟ�ϾQ��%�P�^z'm�i��^�zt���G��i׿�7_Psf-.~�l}��4��2�G�g{�Kc���h���/�k+� ~;FE��S��ϡ鵍�њ])�nk�Z�3�?�a/��� ?��r��A�+ �!�556��+'g��T��-~���s:)++�����%�;���1�]�#�u�zrkd���Z���_&����Y"zAɓ��0q�m��E�v���P9z���t����z~�3��Sn�v�E��`��t?�R�S�9�\�PK&�%%��I������$���=��嘘<J�Q(�z�$�<k��rHN�h����
�������*��i�-�%�c7�^^ƀ�ë��� U���hm/peI=��
''�Tn���9y'�,�a&�0�AU=�b�����zw���|���\�t��7�Z���"Ǹ�^d��u>���?���p��9󃠤�ht}���ŭ� 2P�T�B�aP1:�S"@۠n���5/릅rD#^Sa�����J��ċ����tGC����ń%�Zg7!���m������2M�F�"S�z��:5��7��ǽm�NiF#����m&e�F-o-��qu}�Wx���M_vrHH�1�y bҭٞB=�����b��.ڌ�cړt3_+�}N�hEhY�h�$�W*��g��:|��k���^j�8��c���0�/��'p��M��C3�!S�+��J�#�(�zkG1�Q�xB��Hm�E�khIO�c�-�R���լf���m�\����>��s=]��'����`��U;U����ή?�~i���(L7���|1 ;�^/��E�g�p�O��8o꨺�X(Y����*�� P�?�z���E�V�҂��L����>u��։(����%%+#c���!����os��KaG$
;����u�M�����ɒ�@*S��c�˘�i��^��mtW���8�~Kq=*)�$r�$q���F�,�<Qm��O�D����O� ��0Κ{P7e9:2b�~��S�h/�¾a<�4�(��U�fRƙ|OA�cS7r��+Xu��R>��B1�4~h(㏊�yyRrF���0~RX��c�L�(<D����ol��6�½۱��&U����G�����:�	i�P�n`�����W��Z�0w�ɕ�R0������ԋ��vӁI�)Uf$��x����L�d��h�=��	��ѥ��K�����k|B�n���Im���+�H�9ئ1p�o~P�rG����F����B#�\0Kv@��f|(��Uǵ�H:!��{��2���ɪ�|�SA����}�2r��-��i�B�_
e��T<%t.R#�_��%Y�I��u��PZ�%�� ����=��t�?�n�j��s!��J��Ǭa�j0|@����<�=�3ك���r���ɩ��a���<P��q��-+�[;����h����
��t�����j���^"�PR�d���diZ���O^��L�z�^NXޞ�5>>Um��M�b&�U/�gB�v�׈������u�p��X����<�X�4IrW�bb���J����T75	f��x����53�B��h�c+�N{���cC���-��ص�\&_�9²Z3N�1��~��A�N�ӧO./4��9���cc9��v3߅�J�o�N7���re�|�t�u7�um����8��:z��[K�<wI���e���K��rD��fv�Y�03�:�b��SP���'���u�iG��= �G�~A���8Ƿj�CuTU��'���m�N&ܟX��Z9v�с$):3��d�s�6��$I#?�?��]�>���ߨL�Wײ�S+|�n�۵D;3<e	�8=���GDBͫ�nE*�c"w~f���lT���}]��D��4G���+�uf�6��:�������.d�����j[���;������c>���,.fAe$Ń�����6ϔ(�ʥx<�?vs������,	 6 �R�g��B�?�J��m;J�j����ōG��FUm��]dx�8��W������f
�V��P�w��u�b�qGP�7�=<�+T��H��ίG�'FB�b�ފ�ۚ�M��f(!Ǳ�?��쥤��U[�^h(V_�G�G% �?9y~II5o�>�J&W�<[�ccc���ܙIN���nz}��n������/៊���(��,%.�%�P�}�P[{�f�A��_����RRW�մ������4�x����p��~}���Ծ�Nz�[��e���=$or�Z��N&'[�Xh6�L�!��D.sd 
.�&��*�)ccE�����F��~4�e,}�x�\�20�t��B�f�<'���G�>{�5�ړ=h(N8B�ɸ��'᨞��V'�!�[�����R�Jt���/�r2�+�����&�<�)��D��|0]4 gjT�ֶ$�����Y�0_]�3��$��$�?��Т���- ��@}�F�u-�-vF��ʚ�n*݋o6��U�O��p��%Ѫ�Z92�{��'��-�^?�Ǎ0}64Ð��˜���2\�;�?p���"�-�&&&,���J�װ�]p���J���>���A�Z���S1��R��Me�館4������ 5�#ZK�߳�{��� O����t3Z���`����ju�8�����q`�;�.+�Nr9`�����r�0"]��!��y:mҒ���BA}�q(�̿h�D���~�}=��Uo������E�Lj�K0�2�{0'�1
�G6�e�a�b��n%�^W.��=HLNN޿��w���y.��\��-%ؙ���:c2T�4�~���`����u���(-gy��Hz8��r}��(^$��c�d�l|����oky�VW8/�o���~JA��^�\> Y�
֒��v�ڑC{_�5�rٿJެ�e���&�u�V9n�����v�ceu5�c�%e�����ˣ	�y��A/P��Ō�#?��hN��G�;sGm���� !�}S����������saBN��<d�Q���{�o�A`j�~��h���B@@`}s�w<R�(NR��w�����xy�9�M��#hj2W�����{�{���?��) ��~����a?-ud5x�o��3Ivǹ���K��5fe�0��)Ǥ�B��A�	l�Cm]��f��oB����S�Ǹ������g+P9uo����ļmq�=5���޲㌣?J�>�%%�P��d�3`m�&�S��5{�����V��"A�vU*jk?���J"NEB�~12hu`DTY=���F��CRN��eC�&�$Y�S���mm�����=X8��<�0�3W���X�
>_�ݳ�s[,�w
��@0������ث�e��v}(r> ӳݎ�� ����F��2�r����P�����&SC�}y3jy4�h�~f�'>ઈ��ENC~�TF�2�r�]�����ӽt
�C��p2n�Z����@�ä��$���UϷ]#�{6��Z-�p��+��KX6�	�	�p୭H-�_Y�f�:��a�J�d������?磀'���D�����T	#�������8-�J�:m��:N׶���܁����W�U�i�e��E���:M����?���*���!��V�I=���VvSSh+�Ϯ��	0�H�S���{���9���SQ]�e)z�0��5���lg�ˉ���	2��6Mu怭6�E2��4��c�BJ^�~�a��f�Roj�aKޠ��*��/���M������,��x!����9�{~�� ���p\�WݬJ�Z�x�f����É�LQ��kd�3�71�����K�l�N��P�BhGF��X�\ҋ�~'б��2��EB��_r|E�Y�W��#�0�����^Aq]~��5�d�hǧGT)��m��������s&1lx���<�d6ڐi��h�t[��C6 ����	k�|4,c����+	7'��x47j-�y
n���8�"t�%��0���
,���Z�L�X��vz��u(���\���q���g{ˀQ�*=����������^2��5������sv�k�ܶ�]��ܯ����зڷ�;���&����!���ʑ����Gl����ʰ�k�\B�%��y��+�jj�P�R�rM�l{8ƣ��5��~����]��|���v~�n9�k`T�����`�}���*�O%q�(�.�z���ߟ�O�1�e�u?�
�ݩ���� \��b����`3�l^圈؈�%�W�t�_?�d�>�w��������h��s�-�ɼ����	�P���s�ig
�=��ˤ�(��S�'���l�Ar��7r^�l7����ѽEù�	Y�;ѿ��BP��HND?�n�y�ɮa���X,����Ƴ�	b�VvY��ᢹ`\U���o��'�k*'_�ɗ���H4�9y�wY��r���K�u��Db�zX������ݻ�h����&������[��:Y�e�D`_�b��M�K�0����_ǋ��L�
HH�w����"��:osLY��/쏞$#܈HJ��3�<�z(T�5DL��Ie[x�v�&�x2�8���s��J���yyP��z � S-}�I��EI�U�e���{[�:+�׆��V��W���&��,Yw*W�ṠJÓG?�h#�ĕ��A�r�&\�d�dڪ������ o6K��~6���K+�$�P�[��W���<1����X �K�o�w��*���*v�����8�S�(ZJ��Cq8��o��~!}��H����-�Fhn��֣1E��G̓OdP.[��Ժ������������}N����ꂪ*��q�Յ 	%��rF%�`]t��蔡�ў��J �?+EQH�%w�L�q�'�)�9�%M�Q��d]B�8�:�9l�uY�:���o9iV�a�3�T7!>��&G���g�j���(�9`k�?@��%)o_���=�NV��s�o�|K }�,�`C����lc���x@�C�h<׿�˅M"�l�z�2ɹ������)K�u�76~�҈�kT`A[��&��[[}�ǡ��>^O��'(�eߣC�eX1��w�7ӣ?%IRyw�?��%��sQ7�Q$�ht�Ӵ<>����#�����]��p�n>�����"��vގ�n�ԍ?<-�����̫���":D��F�4�����J@T�$�)����"i���%�L���$O/���ᛤ	ֲ���._��n����Q�%ȷ�����]�~��b����_��ղ�e-I��t��,��~�9�W,u.�{�9'�\O��>̷I��?��ke��}u���_j<H�qT�6
��>�C����^'萴K�a��0O�Ϋmń<�9�H
�4�zU�ʶ�J�����H�y41������)/���6���o�N]/��h�8�B��9^}m�a_2x�F��N�
)w�pdQQQ���������
�\Ff2~>n&v�I��a�C�=[u�7�3��Qo/�	��]��?|�-�cX>n�U�1�c wL�TXc^c����X5V [?��	����\�,VɌO4ҫ��h:���3��C��
&�F_6�����O��0(�g���H�ݮo����ڴNz�<֯WbCJsr�}���/�����@���+{��n�.�:(�	�M�~#QQ�9����ϧ�$��V����x�g�E�^[��M�<)r�?(�wZ0{�s`�G�PcyW��	`����.n+2��C���$i�w�r�D��7���3���#6v�<,%�z%bz�ֹz>�ny	�%OM�1ߵ���J��X�᷑��y�d���i7J�J"�8r�(A�e%z�� �t�t��c��dq!&�BͅQ3��������Q���YIcU��|�H����e�Rc�ӗ�'n;*�/�G��Γa��k��-�:VV�/]����)�$���������j�c(�j{�z�g[?�_XX�������I�ˍ����,\^6�I��{]�U����h�d�3�%A���U+����c.���k�%�����^#�̗L��]
X:%P/�u�G�?\�ݵn{]K���s�c��{̲φ�E���.�����;X(�Z:D�=��3��I�L�r��]ԥ��Pߛh��ҔV.y��q�:���ڭt[
i?�
�W~v�; n��)ϫj�%�ĉ���I���$/�5�'������n����m�F{��POBuu�Yk|� Ql������W��Q���i����t�c�H�F�J��;��$K�!�"�EJ��妛[ x�ё#X�Xg�b����Ԕ��qx_��V�"������K�SҰ���F$=j�qY�NfQ����� ��8-��;��[0�-�l��,�R��̲L�@��>j�R���c?*mQ���#p�߯AϞ0��H\Y�k���_4=0�@t
�z�M�px��^y:Qux'�La���{�8Tj#�\D9B�耹�98�l��q([	�~������c
��FEk�~�Bc�^9���>��i�,� u�}�����A��ô�Z�q�{
9@�fB�+�b�-{��n��`2�?�K��S^����H�9�	��`�]@$�p��p�T��t[�$�Q2[�٩�`�B��
m�#�t}�<��/��o�5�X����a�s)?�i�
����g���2{�i��zT?���08����d��y-�ԋG���@.���u��,sG�a�G�������V���:~�1������X����e`��<��	���@3��R�յr �y/��y�XHb"QeE��� �0�rG�$�ϭv���Y�|`������TfNw�r'����,��G��Ρ���MW2Rr�����G�u��l_����j1���e�Z��T]����t>z^T�0Tqh^T[�3))	#Y�H:w�W�A���Lɯ_���E�������#^�X������ⲥ��Cs��7�`����$�/q���غ+���Y�qε�J�,ĺ��q0;N��y���`�� �}��S/�`�K��U)��+�i�׭��l�9��5EO�d����W�<�{�zu��n'���A�Ļ��]�I>���>�ʵ��"w���B��b�o	ah)�YAhKM�H�PV��u"����"2rl�vC��X�w	��/���qh(��ȓO!!8���sAt�za9V�I�!�i��6����Nua=۩gy�~������'�ڞ1�,��X���1$���!��uo6Ԛ�b֭E��y��҆Vل�at(���朣Sj�;ZFE�{M��.%�H�<i��{�S��<R�ؔM��]q��\�E�\ta�_B�/�\�-O:�F�-\^��kYzU�[lI� �7|-�iZ����RdT�4j����	ͯzyU��J^)� L#+SSZ�����\I�Ѡ�^���ia�/9'+k��?*��xsr�9_��H.��x6/� C�g	9߇�Hc�8i�� F&3�}\˳��2���t��ȋX���l�d�I��e��ȝ�-����PH>;�nf8`�M��M�eΜ|���?��`8^۴�Q�Ӕ�CH� ���p��I�����v�����E���eSy��us'�	lfp�ɣ����y2G��J���_�����6�FF�
v��Sሂb� ���am�4�V�Ы��C#��^,��D2�]�A�<,��&��x:Τ_^�a�k��]�4����\�2���ܴ�Y��?��o8:��04�������*?|^�Ѻ��:e�,�,���r ���T_@D!��,@�G%����]6AB�3`c�ZO-�#08��,:�#������c�T�.����Z<���s��kC����֥PCi U��-�^�;�B��b�����e�ٸ�'�Q����]��6[��Q��,ź����6d�W�3F�T]���]���ְ��̏��6*N�fT��5H�
~�Y�[��W�L�\��
"&�b&`�v���^^�o4���(��߿�u��907�����W�(������
�ngg��6�c߿pL+�NN��-;�6K�J.b�eK�>'��G߮���o�u��[��^���6�=+�������<�^|)���j?�N��9D��a��-��������zi�1xy�d�Gɱ��Q��lV��ٖ����ؚ�~y�z�P�9����Pd���Cd�k��W��l��T�K�8�x�m�&�9�p���A;��*^��,��ҲX�$���>Ȅz8�0�ٖ2-e��RA�A��]+c�5ȥ����$y�L�iK���(X3��L�(>�`�h����~���)y��EEE�Ke�*i���+"22��v2�ttV�2�q<Uw�k�U��X9�{W��C���5�$���Jt��s�c��梯;4�c�.�����仜w��J��~[o�2�Rf�~|i���u�{�4�-���U��q�w�{֟��h��(4B�T��0TA��^)�k0�};��]��3���y��C,��m�삂�t%J\��m|���Rmm�֏�]�fݪ4��پ�(T���5���YR���ln7/_�s��y:
��*&X�\��j&�HF!��+�؜�r��`(���ϩ:\��ٝS��C%�y.+.�U�m����.��Q��A�/C�c���D���ySc7�s{�KW���!����ŏ!�ێ��N]{O��t p��zF�B�H>��3�׾a���m���;a'f�yď��X���1G�r�ix(Ǒb�$�����Fm'�S�U�\���&��WWÇ�z]'�~��Bk��|�)���p8���c�A��;��y����������ߟ���:7ȱ=x��wc��;J�0��q6/��QX�f�.���U�L�y^�7+$e;2��G�[@Eټq�4H� ���tw(H7H�K�tHwK�"�t�"�"���]�����Ι{8gٝ�����uϘɶ�E���\{�}�7�4Y���o�o�;�9��]���Gy� �B��ɭ�i�� p:	�G��Ղ��L	]�csu����MM�"�����\��^�Wb0���Ƨ)�Z�P��|g��x��o�F�9�,V�ڑ�����{��ԯ|��S<��orF{����A�+��^���SMM��S:B��)��px�M�*X���Z�TdR�����I8�kR�rL$�'j:��U+K��e�d|�}{��2,i��÷o�*�5�x򦿫6y���:\��uQ%��=��OÆ�5��]O]�����T++�U������]������UW��zZ��B ��ϗ����"c����Zb��ML�0��⣣�_��LxR�O���в�7e)�����r;$�Ǌ&�����i�2=+>֞:9;������#Z���  \�d��'�n�����u+�����N����G)����������z�����P�u{�<e�9�Q���NMܼn�R��m+M��M��a���"n�z��x��Fa��F,ӂ�����D��M���#�Oƪ�E>�F9����4�j��Q&�u�Tk&�ͫئ����T�N���Vk=Ѱ_RR�jP³L<L�ə�"={�E �K�{�"0a�=���n�5`�LMԎ}����2=�~��@F���x ��\ӵ׵�w��ATE��� �%�Fֈ{�B)�?W*;���K�V���/�6��M����SN.ZԿ(t֦�L��]�E8s�[�iH����]b{�kH2:
�m$��I�foZUJ�h�Ij���G3����K��M5�Q��yٲ� �Ju��e4[���",#J�x���vc1{@�6�ʜܲ� �;���-��{f�-R¥�[/�L�]d����|���[�:����02�Ҥ߼W�r~��[����U f�
1z����F_�֫!�=J�-=!G��u����Ϻ&�	ϯ���TÉ��'��!OW[���}p�A� ��	䲠�M����c\B��ť�����a��z�7�3�[qC�/�D��R(�x�:�$s����tx�Ջ}�(d�B��d���q���8���ʭe�������u�v]]lS�m&7<���W@I5ߟ��W�'��Σz(z<eR-�|����)��\�<��������������ޮ(o���[�)u���cqy{�����=t���l��9$0����5��WR��3G~S���Ho�{�LpK�b��Ȩ:z�~9cE����*���ɿU��Ըc�Z����7SJs�_�GӢ6��n,�O��!�N#�ɘ�.�!�e��?[4$���9;]����M!x��~��X�Os��`�5F>�Kz��'�e�^Ђ�Tc����x���Oy���mf�S�2��ܟԒ�����3�4@�Gɱ[�$f���ϒ��ۂ
��"��[-\	���\�~Ϯx�R][����o_�� +r���1��_���*;��la����{Gr#[�Q"�����vѥ��h6�����#|w���"'ǲW��,������ �Xd�V&&�kڟ>�e*�V��������K��J��XM�yg�ۨ|������B�Q����Յ����~WW�f�x��/R�gL�lYF�X���'�'E�p=�*�W>c���fs�{�&#?��$Q��N�Z~嫝���N����k�֐︕z����T�8LhV˲a��]�_
k%�vB�Uz��
:���,p+7J|sx��t�� �ַ�1/�sǽP���sU��������[��O�j��_I���]a��=Le}�gN�?L�T+RCdrg�y�������_��Ԓ�H����VT(�
�E�ک���lq� 	1���ַ���w]t�V�!E���p���8d�~���������Q�:�<�l�����enn���"U���z�!:&f��[Hy9��V�X���d��(((t@��c�~�����p7��a%��Z�MS8ꦭ���z��H���:4�imS���W�o@��0�}�qwuq�N��O��	*���i�
X��+a�	�1C�.f�3�,����?��ba��L�]��T�z^�Z�����"*� p�{j*��@��T�5><�Z�0��q�( �
��^�}�����w��4��-n[������xDRo�\���|��*S��L� �9<��e�X��s֢Y#G2�]"�R����f�k�z��ב6�Z�Q^P��I����װg<c(E<��f� ���]�����f�8�k{�B5��>�j_��vfQ�@u �,L�a�'Kv/R���p���q�HYۮ���ͥ0����7�ګ���LݎV|�{�;T*99�x
���i>�!s��H%�~(��iJ�/<k�V�e����MX��.r9���G����֮D�_��͵��+m���A��&��k7�M�벏�B�� �ʣȷ��DO�{�U��	n�׎�ɝ�l�ií5��,~|Vũp���ם$�����������[WL���_k���L͵[��O[l5�2�Gs܊�����S*@\v��ŴQ�D��Q9��,]ڈ�F�����xȥ���K�l�Ҩ�����G8�1:?~`o�w2<�?�{��W���N�ͶKۑ��N�Q�1��7�3't��^S0�Y�
��[��-��ބ����"��f����i�QJa>�h��P���I����v1gљťҵ�G��1�����?<E���$x��}N�-dn��'Уۻ煌�m�~��?����΀��u�~�������l�h���K,��`X}.&!E}Gd|�Z22���O�>w��#�Sg�Oj��l�Tppu\/��^���\�q|�z�^�$j��sI�O8��ށ�Nv�tb�<�O+�u�6�+�.���>���?�lM�\vJT0���Kl��mg<%yS�TaV���w���@���ˁ�ҵpip�; �?owkhY�bf��kh���N�Rl`)Y�i*����eo~^���GŌ� ��E^,�UU-�Ga�ށH��%��t�b#���U�����{#Y+I>�֤]ta%�T���9�tr#���3e�D���Z~C`3X^ET����a��F�:���� ���zd7<����6���ԛa*m��k�|�Uz�Ӽӂ�|!�A������YvwZ$�uw��L�C��yC�ի���k2���=��i��m�͙t��3��;K7#�N:[,MC\�؇\�d�j��/Hd�>.T��^���f��Ȩb``���������0`�c���@`=�>^V��y>�-�\0�-�)ɲ�I0��9��$-$��ejxz�_�����w;�c1aG:l�zT�?�����-?����S�S�xΩ�Kn�(����y}�¼�:��{�gHhf���:&�
|J�釣,�FN���CL�ﶆƇ��*R��nw�۪���r��]�BԊ1�2���A��?�*uO_��L�_�2���a��lU�ҟݒ;���k��u~�ʪ��a��ɗO�Ƌ��(Q("��_��n�H�P���lL0���,rA@�8�2�P�7ӰcN�RM&
k���.w��Jc5b �Յi0�K��v�e��0y��"z�ud�8͇��>�]e8��T���=�;obf�$�R7x����c;EMd�C�q�T�v�Hz�,��X���p�ZׂR�����)C�n����բ�֬3�j���Y�w��^���T�l���'w�t�����ǵ쯇j(e~{��im��+���@h��/3T�IIH��z�"N��U�9'�KS7Q�Z8�<�^�
�յٳG�|Zy�f�4��z���!�s�`�w=b;E�-���?�8J���������kz�д��[��A������piH}�t�3~������	��5>O�^u:O��]�Fx���U��$b�,3YJ�,�_��[:�ߣ��ݮ���R�k�A
�ܭ�eCp^8	}N�������MMX�Iz?a<	mK����+�-�t�r�%I$P��2q��ڡ^af��$1��L9$�K�N�5 �9U�VeU�m��O<�����o��a�
P9ac��{�~`"U�R署��0!h~qR"��#�~����V�.S�\�r����b����O��%1�@�oUUx���"W��U �,��=GG	j��yk�qMމQ��9E��k$3--�?��{	�E�h���i��$G���� =Y�)sp�}�H�����x�]���K9���q$�߽�����GO��M��JkR~b�}���i���t� �V��̘%���?��6$>�D��6�������j�� r؟y�� 2�#�*"P�9���G��v+��B��؇Ł OU��(����N���c�Z��*����P,�="_>>�f�;�8^K�?���]&2���0���NQZDo�z�N}4z|���;��$�j]�S��~Z�MO~o�j��q=�Š%e�.v�X���0��~������,#�.i�/�*]rK�Y�Zy�G��}=��cf�7�o���А��4*<�c�1^�d� ��wq�k�����+ה�qg�Z^�YQZc
p�'�d�
�hQ����ػ mˆ@fj,qΙ�7/<i��-E9G�:�c�?�)��÷�a:ޘN�١�\��g���=h��f�قV
�>ڃx�h;|n�S+XlA�M�qT�M�����ݑ��W���i��18p�Ә���͘j�[z���e�?�|�cy��j��Q�uj����WF����ă�@�,0���&���S1-�Ϻ��{���a�O�����!�h9ҿ�Z)��ـ'*�����4dv���k���h	��x�e�Ǚv�n��n=2&������A��f-���~[�\���d����?�[�߄�#fe�R�������-h;Ƚ�o��/A���"��~p'L �fL��&�H���@����gv�*����CP��/ם��>/8tam�7gZs��	猦ډg2}�R�@����/����p��(1lj���}�Դ�F�Wh�M�P?�Xy296j�!;6�h�A����U�n�Ջc�FG����|�wf����5Ͷ�ca��n�>.҄^������7�6���Է��Än���j��]�FM�6�X�:Ժ�s�A�Q#zBBC��
�`Q��D�jX��[8�kM*++� ������P ���W�lZNEOxB���(�Q	��;�t7�sR�2k.�Ӯ폂܊\�35�A�[]i\���5�~ch�J�h��̠��D;GqѨ��A�N�Nw�c�zSPh��d]�t��O�Oǹ+VX�m�>�����a�铻/
��؄�?��B�H�3^5s���q+,zW�a.cڤ�]�>�Ƙ�n�鹈�H��tQ�O�7Ci\�|�.�IIIK�zqey鳙V���ҸHh&��V��@"���愤�������N<��5���ɒ�'�o��f�@CB &&���I� _�;�Ķ�嬤�X�2vG�/���E���3y��.[ޗ��/�ڒ���,:�S����`>\�,e�~��aa�l�X�~%��Ĳ�H���ܮ�=��vz�N�VVV������K�g�ܼ��>D N-δ/]�)�zcK�z|5�$�G-jdL�����H�e_���E��#|h:<��O�:��Z&����j[��[��8^����E����,�Ê��[Ea8lW����k1�X��h�󛶥�M^�[���#��:�g�Z/����7���޴�Tk>-��������T�>�r���}�%�_�\�Ч��r�LI�_=>>ZS��������c���28�g�Ib�Ј�Z����\�����,�����v6o��L��bF�d�Fv����j̜�k"O���z��q���Y��@"#o<����C��yy��{{M���KQ��^���{	3��m^�f6�$�u�*O�ﾚ�(���o�g�T��M@�s� �E�������8g`�݊_tz��R7���J��OJ�+���a�9�������U�&��ƭo�h"�Hj\�94���"�هP�X�#��^TTG���:;]Q\�������$��J-i�W���݋P*��{p =`�T���gu�������~t��:�7��Gz<�NB���cY�.����w�rvWlEֶ��Tf�lw���J����~+-!e�sVl\�FĔ��M��z�Lm%]����^�YLU�%�e�e)@!!�.�lV���9�]`��+���y�y�j��_��=j�뽠���e���xx�E��|�y��x�������j�K�����$�,���"���O�v(k2���ۈӈt����<|�r�� ƺ��B�2��G~,��|�v4���$�0oߎ%��)�!{��_%@G�w��(p)�5�H>�����O�~��U�����:ɿ����؃�8�bw��R��]�=Q@�N�?��S�J{_�%,�{�yOƫ$ؐkK"\R.y��R�x�6O��>�.t�H%�5d�ϡQ=�ss��%�><iu�}����YJ�����`��r�y��O�tJ$�v�r��8�,���6�WȠ��w[�6�7��6������#:�`q]`�ND3��e SWͶM/�W�h"x�U��$ �n0]�����������+g7��/J���j�"��>0��pĽx��ɋ�`���0K\\ ��Hj�����'4����|�g��ʚ~rlaJrQob�		)eOA[��xvd͐^������6�6�O^k_$Z���-jv�ʹ%�4lĴ`�5�{���?��tMeEK�PD>=f����c�<��2` ��8c�r��'�.'���#g)�����Y����F)ܱ�&t^��]��0څ�)	��b34}����.����gb����`�P�/��D�����7n����P�@I����Ns���e�؇u��W��\cI�~3d/�����Z-D���@�¼X��T�#��#YB��?�Kh��.p����nE�f�M�"R~�-��P�Yt�)*�[G��:�R~�	-���[#A~u����̜�6�:�����T~�$);w��p춠��X�˪�I�TK�9������g�qW)�{�K^�%QϮzc�)����w�Oʘ�$	���	�q��桡ܸ��^DˎON+f�v��޿K0��*V?	��ڞ�.:�2����:Rs�:,�,����B�3P�]iiSS��n�ᦽ1�J%��u�z:��N��퍕��R�?L�=�_D�+��a��~�zS����KR1{:���[ڴJ�y�9���BD�pp��%^ԑ���Ͷ�����!7��l�x�t7A������?��ц_��L���(���%��-����������lU;:����7�BJM����hU��޵cOh# \ �|Ê��w��'��Q��Nҁ�KYB�i��a�^���fl_�����^BCC*VG���� ?��E��T����B9�M��]��~J�������{�n�bu��f#����Z��o��|�t��$x��왽=�m9>U'�Ѿ^�j��4-�U�����^����nl��<�U��rd���.�}V�Wy���&9k���K�+K����Q��&�'�����gK�?n�q����@$x�a�g��?h�������qI7+B�J*�Gk��>�E��<Z���F���.B7�$�9p[�X�v�	?��^�Q�򥣴n��G\��Y��;T�6Cć	�kS�Vچt�A���L�K���G� �kC=y�Ҕ�&�#^��KI!��9o<髠�Ɍ}4�]��7n62�Y��~��2S���n�y./|� �1`ط"&܍b~�7�i��D���c���%�����e�غ8?/�9����<S�t�R�j!e��'�#�
ITS�L݉��Z^�I�S�'�7��Ȼ��"I��5�
�ف��E'j���u��c�	c�t�����&�ol�� �@N#c��LB\3T��|����D�����A�(�7l�x1�յ�2�f��Nh���ZP�^�5�U-�ʞ����y�k�*;B���NGS�
�Ю1W��h}6�i�i�ơ��6t@X�>�Up`e;Uک��	�F�N�[1l�O��O�l�{b��;�tB荈�gr���}?��Ղ�K��):k��4��E����O��b�",�s�)<Ї��^!d���=�Y�P�c�v�)E�.�q�Q�>�]�������jJ?0�3�+I�Z˽�I-Y���ngx�@���g�"��dW�Q��5(n���A�o�d��(C��_/�Og�dg"#�Ƅ4��<�i<�ͥ��j�Z��	�Hq[�ϊƻ�]!D&���d'9�����e{�مմS<�e���<i���ߠs������D߼��_8�>w�49�����gU�-�L+���F����<I�Tǧ��@�y������Y�A��,�~�^����M�vf~n����z��-�w|C�˽M
yG�ߍW�`���8��C��gf~kߝ�ZeA@����
+PV!��O�q�_��ު>�u��X���g:�����y]ϚB��D���-.t;g"�-���!bf��m:N�B�j�mצ���L���Y���5]�n�'�8ł
�g��f�gp>>>ڵV���ŏ?�kL��y ��G<���cD��Di�s��*�Ol�ZԯO�,)Ը6Q�U{W*	���)��`��*;�s0��W.<���aV-((p��ۻ��7_#[/q9�Y3�YH�SaJc����Y�怨X:��)i�
�Ɔ��>�pL��ts=��sJ��gCv���j"��({ݻ�~h��{�}iHqsy�>������nV��~��+��{T�a_̆�x�JӮf�_���,�}!�)�R�h�7H��V�6�7#�<PX�kC.d���[JV"i�*�~�☥-d�R�oޠ�X���(�u�,[� Mb�JH�ݽarcH^Q�G�7y�S��;�Ʉ���g>�$��r�)�+�|"�1�3e����(?��Y�{�??�I��[��F�r4�; u`���A�0p�F�&�fJ�l�6 �g���u��~�mO{�Qa�S��D�~���]t�cZ��c���I<�w�@�nP�����+NrZc>�nP����r�=�x��I�=��j=�u�xSY�;���>�X<*� &B�p�y��.�Vр��7I��&����8��(Q}� ���v����t ��:��h��N� ���(��I�bfA#��j�'7�P���N��D�[ ���� C�y�q�Ix�Ȑ�xJnR>! �śڳ�ꌿL/�I{o�p{�в���e���0�v���Ne���1$��*��)�^w�N_�Rs7�E��>��o85:���~?T�ڿ�S"���ykDFK+u�\噖���J�O	������5��u|D��W����@W�|����~S+�V�_M��?�i���R]�;z�\�^��N�^�q�K"��r�tΧ����	��lX�їH�]�{���L��@�7��w���nݳL+��l|>�*d><,*�}ቶ`ta�����[C��I<�w	���5Xc<���<�_�%F-sm�-P����% �8��p�;yR��`�j>��Ɯ6O��8�j<�f	q�A���ay!��E�9�e����PM-1w+?I��������s�Ol�Զ�/�m���{<��P��O��	q�H����;Us^^���+M[�R�?�_ӜN��V�;��m8����f��ַ�1�ϓ���~}*|r>�O:dZY�~Hܘ>>2͟��5G^��v��#9��Ϛ������'��$�Ԙ�,JG-�m�a�~�^�����2�݃e�as4gPL�5)�bҷu�*ޢ�m�����>CF�s�ξ�
N:�qQ�n5����-��`K�b�	�r(����	�Ҕ��t���"���7�&�7~#��a֎i��*SX%���� 5]d�F�9Z��v���D�?�9����Dx%�����gw��f�R��2`�\�О�B��Iǎ���H{wtE�7l��^@�n}�S���������LK^�ʝ��)����P����䙻��8m�F!%Y�����0����eՍ�U���\�?^���F�YQR�kK���q�A�H���d@g�z��z�H�h�h:1FI3G�+X����
t�h{6�b�F�����sw{t�+Xhd�v�Ш�}�p�+��UڥV�}��z�ۂ�o1���ʥ�B�{�U�4�G��95釸](1$��w�Ì<g�]��nI����b��f���f���p�mX���F$Ϳ`Sy�����t[�p�40dM���J�E"��Wz	E������\�o�Nə�g,>Sd:y)�(���VO�b~��{��Phx㘀�T=�v%\�fُ������͝�5)<�Ir��+薴����!]CP(􅺔�+ŉ�`*{oO4	(���]�P6́F������u.8�����F9��/zȀ��g����p5�l�&����pɪ�%��4d�>lUP���,�w��<�|��Gr��b@:���\�ݑ��Q*��}��@��ޙ�m��9�;
�<����\�k��W�<���iZ+�ʦF���cLI5=ފM��N��=�<�Uo
n�K~\�H|MQ���P'��x)�؞�QyC����,�ט����w�������c���<iJk8�X�K.�[q��O����*𽈎��JU��m�,9���˻�>�byY�0�N��	-�3�����|��cV,T4�{���n���Л�خU��Վx:�8��J�n���ZmM�g��V����|�~^�2��ꯊ�����W.�A"�aq��q"43�eq����}b��zk�Ǭ�߯�����A����Wwm�#�1u�N��>�㋓�y�k�_��|�[~�-�9p��'���mA������Kt�lE����)h����S��V�Z=�^7�Ӡ!S�������TŒl_x�24f�L��\}�� .�#'�%4�dI�/8���d��@|/Xu��gl]ڽ"���Ɖ���;��p���s��R-�J����&�缾�wS�
W��e6J�������=�w����hk�?S�*�k�]�Z2�pK������-�ul8����Ƌs���{��T�t]������o��Z�긚�'�����,�i
Ps�e�.b�doN�m��SZ5�d�O�0��%�!�>��eR�dlv����mB������M�qL�ܿ�,�7</���Лp�}�N���8�\,z~t���e��yߚ�4G6^�"�[�'�ָF n���hk
9͎R�~'�����Ŷ�u��%�������)M �����d��-�\jqS����T���+R6�&Yn��1����L�l�}l�
�l������ߘ��������>�.�o��Ã�}uxx
p�v{����`;���%qKZb�����e�@�;�R鶾�>n8 P�ʻ8�����D��m�//I�X �* q���o']�٥x�|���B�
 �H�ɗ���X�6����e}��]�3˰'��Ӗ��ΩBE8�F�_�(�M�ce�U9��#�����7�'S��ˏ(.|l|(c.ge�e�Pl:/�4�2���xb�K&]1ݥh���{%�����Em}Ո��}3�RlZp�J|*����Cii==�͡����zG�˔�����L��a^�;i�^�8zy�OO�.-�_]�>�[��~��̽��H�@���(��U��mԠ8.���~�g��-�;g�=�W���9�]�-��:j�h�I����m� #���c?��nK�\�N��<�'l4���ID������ܒ�b[��!�1}n�ٕ\��	8��n	�>���\��lo�,��A���E������� ڧ֖�^5��9�������OQ���}á�%����c3r�x�U�In���s[Qz�w0Y}q�碴Y�����/|4��������R،�h4�=@�a�n����U,�h�ۏ�����~[j����2x�F�Tvn�M�v��D{��"����DK�AC|8YYY���?�S���?�˞)¬�f�@`���^ 1����S�mlG$����)�>�(�F�W/�>
�[V%��@����h�s!��ᇯ��'�a$G,6�Q\Xh��aśhN���"adD$Q���N��3U޾UJZ��Z�,��R`{�V�^^N�@��������;;׬��abaFcac�.y'�h5�L���c���:bu�c�Mx�����~�IC;K�r[t9�J���(`��+�S��@��i���skc��Fv���}g�~�JD�u�%���'��F����.5-Ĳ�KLCy�u3[*�'	v�x"k'd��%Q�jӠ4�j��O�q��
f_�[f��D8d�?b�3u��\1�Qn���$�r��Fy�}w�i�(���8���y��D�'�\� �\���\J|�L		�g�T��:Y[��	u�A�����斖*�Uɡ1*����&�b��Oo��]:�,�����擲���L'H���EP�"�ot�5#=�����Ԩ�׎0�0$��dQ��ȓ��<W������x\ny�8l�&�hdv+����Dc�r�e�
��L:���5:����yyd���	�b�������q�<�A	A��o�G:�W�2�d4E^�7p�ʴ�nT������٥c;/����"��]54��ꁎ�/��/h\�%�s�����?�W?0�i�U���	�0��8Գ�34~Ƚ�� $f�?����c_��V\��Ǎ��N������ �f[�L����m�6)e�����]&گ ���-u�dK�.����_,������Y�칏�-������T�f~@�K�-���c��%x�f�!�e�<+C-�6Sc�u��)U��t9�t��4����[g7����\�Uh�]ͬ]����k�^�}o�gsqw�ki!�k !;�:���ׁmԄ�P����[��7�ayUUx��O�����&�zc�|����I��ǘ[}m'ݩ��6jt���^:V�4�T� ��0�3��ݧ�u�`��\�h����.MSkA�T" 
�)26��(R��ǈpC("-*�3h����ՙ��l�iqѴ�5.2����s>˷��X�#3��@#N�%I�dJD�+���� �U �>���Y5F�A�SaZ%�h�;D���0��Z�Q�K9u?�k(���ʨ�f��P}v��Q�	k�|�6�������#Z��ؗ�^_���0�����c�F��D�u���xzT�ً����$y�"���7����vU��MNjLaOB ������W�����h�ՙ5�E3�Q
'��v��"-�K�w�ĆS��(`D�'����W`Wm �:�H�,�;�``��Zo.���,K���\�di�d���r � ~�C�nB��nF�sss�l�$�P
8T�Ȟ�,�X���Ԅ��8�K6��Ⱦ6S4����Xu n~�O��rl~rl��?�"'':i�Q��l3�\9g~��+�:XX��0(=\�`�K�q���M�� ^�1}�Z\��
fӄ�P��S�B�.��=���U�8I֒n�r�ґYBo��N��=@e&���i�{.8�Dm��抰E<bF�(���=���䁋n;�Y��-��ba�τ�b�"�h`���w��Ld��֎�F�����-z��l�R�B��I��d�
�Pd���s�ZA!����p={(!���r����ZG �L�=�/�3�7��!!(,��h�J���{�B���ʯ�¤�	�Z/�΅��&O�+g	v��(�w|j*��vJ�@~���J�&�'���FO�n��R���i=�Ȃc���<�iŶ�r��E��� �(\S�R�].���|$�\�����Z�x`>�����E�n	��~�!�d4��|Ohu󇍡&�}�?K�Yf�`ۃR�����	�z�˼ܛu�I&�K�?^~��s�Y{��hmuZ]u�d��VV���C�H�Bn�`*4���¸�D��A� )d-�=��6Q���)<�YK���$��n�YuS����))�1Wg븑��c�L�_kve#�D�Wf�i�g5�p*�˓&j��R��X;.���	߫*[7${k�ٻ4�����2=&��m މ�o'+�&&�v��v�N�u.�qs���ꇣ]�V����0���e��=��b�5���VVLG�4�DsB!���2hUR���ӈ������542_l��������1��l��7�@���R�+�����ʸHܼ��/"����lmaxP�VbӨφ$��h2 c�Ud.��!�?�~�!���78��+KK����1'}�������Ss�S�p7��k`���`)�k�J�;h�(�j�G�x�e����e�X�P�����ѯb��@8��~�0��nBX�$�f���L����O:�m��8�r�$���c*/���o�\#��m�NJ��ֲ�
�������W�·��=Ӝ��1n,DRc2��� �������5d8Ӥ�I��O�вx�	~�!�f`��*�����(��B�P����J�QJr��`#)������|U�Ю����g_Q�*���0��H^{<F ��^��5��f�D,)Np��Ԡ�a����n��W���ë�G�N�P��qݒ�S#�[a-M�J�,��Q��<�v-�O��L1��yv�TXe;��
@-���$��n�*�@���0���`OP��(�/�%��}���F{e��7Y����kҗ�4h���d�8Q�7�����R�����Gc4�υ&ma�\���o�����q���\&X���
�'iӈC��:,,������"�{z�����L�+ƿg�݇�o��L!�~Ǝw����>�4���%ڏ�	-�Iǀ+oQ�˔��#���������&�ca�4y��t���;�?�W~�����?[��u�߹����*����)����̓[�wFp�ӿ��j��=�qT�I�E���k�Y^t%�T�-
�(2���+ݚ��+�f�C���Xx���,����vx�W��Ayzo��O� �%���چ���\����#&R���"�m܁�K;W����]}�9_j>�O���i����
�to�!�:T����IZp�_ǎ߆++6,8�}�;����=�����g�n�#i�}�4�"i!d��|=R���(0��'��TI-q�xؼ�0���Q�z�d.�+�|��c�H��T��!�"êj���#;���W��A^:���e��-��zΙ�	4��i�HII�-��N���8��mf�ˊ��f�xU�?�0z\!2�'�[	x/������{>}r勲6����t�r�{�EFEB�Ks�󬐨�~z� �z�Y�W�ŀ��m?1>nkkK0�J��[��;��Ǯv �Z[�&o�,1-G�5kd��ǋ�{�skn-�p�:O��f׽��m>O�2�~����N���l�=N�4^Aޫo���&	@T�qBP5��`�Oa��0�/Mv�9W���}��>�шh���>��F�!	!���������s�aBP�at̪��ls�e�O���2=�[z�7�T���q�N��Q{�� P�}n��bH$��n9M�ǔ�[L �ۻ;���������7G�/�z/��b�*�)���a݃�W�
��߼�	�O�>m��ue[�C���3���Y�����]\�m��x_0���r�ָ�5�I�,�)bK��0~]"�e�~��5��׿�Ѵf޳�ߋb� �AB����)¢a�W�|(		�]!���t��3�+7�U�!�� Y�.°����S���BjZ��(�7 ��v`Z���V�?I�w��'I��ֈ�=�/�v��K��Gb0�[4�F���t�p%N�kM=t�p̫��Z	\���A��E � >�
z�3����˴R�����&oA*�ccp�X�lw����CU�i
�\i��v��) �=�O��F��19�ϕj�\N��nM�Q��t��|���z��Z آ/�)N~`���J�{l�ɡ����畦�3s��?�|���.�A����-��4��X�Ҧ���v����3�J�a���EM���8���8I+�g��Y��^��N�C]�	���ThJp7�"�\:H��	�ѷ�WU�����w���!��(&&�d�Z��ٹ��˅(�H�܍	�Tcb�I���O
�l�aE�Q�*ue�t��_�X������:z�Zo��m����/�yB�o�I\J����!ʰJ��֒AjYD�����~	܏�`
���Uߐ�Bi�R�&|�6
�"�~׭ؠZ�[�ȧyu[�7��ء[˪� ��L7,S�)�!Lq�,hh�f<�*��.��� ��m6�p��#�D���n��Q9����H0��G��I]LZEZN��fD��8�͖���S�v#�in,�׼��c�@|��a�oĵ�.�kNjf��ΰ�v�А�����l�|^_���u�������ea/�|d_z�̮�*�chW�>���133���o����xc3l�
ņ������͘�e�Y�@��o�yf(��.W�����ʆ�m���j���/��.'p~��[�+��B��L��%�\3z�-�r~�(S���&M7E��[��|�B��?�3����,�����7G���^dN�/}c�3f��Z03���}��u�����v�q3x?��԰�Y�YY0���ͤj&J� ;�2֒�l�p
��Vvv�^vV�!f��)��.���@�<՞y�20 b7��$Z�ʹ��]r[r�[|�#���<�-F���҆�o^4n�Ko��u\��������6�&Y��D��j�J��l�ֶ|ww�֣�Az�*�?����M)<v��g�'��d�}����[D&�F>^^p]!@�o�Л��I�ߺ�� ���%�NK�;׬��E	! ܲWm���
�*����/ݍ" �)� ��"��Ҡ(H]����D��A���;/���1w�q_߻g���ٳg��5�T�g{݈�ϟ��:�Z(��jU�T���)��߂��WJA�0먉83'��'�Odv��u�~���-_V����Q��ܙ3U?�xy�[�
��k7�������!�5���f����Xy����I'E<�WW۽𶴆���G�A��1WWY9��gm�h�:t�����.�"hRFٿs�����ď�f����s�v��)gc�B~�5�eH/��p� �'œ���� z3^��
�h1';��;n=|K!�J���Z��ݧ�5����1�o�S�f��{Wҁ��	a�Q��6��p��m��HM�S]9%%��SV�c��Ʃ�#�h�����z��)�̬���X��q*.�<O�<��������
�a,�0�3�t_�[?�X_j֛��5�g�����K�k��qO44K��$��NE�П��-u�_�D!��[��$�'w��=F��;Ư�F���A�՘ ��	g�IZX�}{֕�ض�� Ha^��X1müX�z}����7s�X3�'O��0��t�^V2���T���MR�O4@�zA����i-�U2������_�9��v�z_s4���Z�^W�	a� ��,.�zJ�Ȼ�)xT��,�J#g(!� � 5��db�>@����, D9I�����O:[��.�n.j.�����*-�uRw��X��p$~��i��$�n����������t��i����	�����.�
Y{�Z~�`k������R�=#����� �ڭ��|�?�1�`����;}�d��St��̳Z$;��t��唜-�����]e:��Ч��ӓ�����[�P1��&�PE�f\Q�e~�l�H����3>�a]e�F$�|�Gq!�y���Ne��bD�j�8�l�$�hW#7:�Gm��Pބ���̵'L/t=�)��;g���>t�})�c�]��E�6"qCΫs�U��ϯ���ï�ő�Y-	�Ǐ>�),��p3����.���ֺ�/}+�!Ұp���B]��x=`	�f�e�	���B�i0��ˀU��9�6_0�v�fg����ؽ�2�VR�-�?�s���i���T��v�}�����Ϳ�B��``���D)�yA��<,_������M�Kꥎ�5�J���=��W�Ax����&�XyKA�qn�o����#��D��j��A�t�j�Yy��c����|��$i�ae�G�� �� ��� t�V~0é�1��tL�'z��H-�F��Uu���΍���~�aאˌ)�Z�+�=��w�ҡuv�qa�]�~ w�7����4�]��V��U�}�I(k�F�����}�uT� �D���=�����ā��^F�3�����8���[��E���Ʊ��tHt�O�~7
^M�!��� ����h�u!�h��P_��:nM�����v��E�W���H`xG�쩻hף�1z�����YYL��+$:X1�t�#+�!]4�g��}[h@��V�g	�h�-֏4�X��z��y��L�PU,!!��֙DPx��
 ���E�Ǻ����!�NNvwS,���?��P�X��-�ڕ~����є�� �[��qzͤ݁�����A@9M)i3�o+��.%%�K8����Bw���ȁdӂm-tJ�)��P]�ǀ��F���Y�	��_�)!G��\�a�-����9k$�zQP�I����@X�`,I�3�w�F<tz����bɨ�QS��Q�\j�ܼ��hR��n~#�p�	Ob�>Q��^��	;�S�0K�S䖎9r��X"!%�뿋��������Puk����`Dp�1�����m��F�4���,?��޻
S�w|�M�`�p�-De��b����%`�^^b`Q|[��O�3��{޹s�t��3�*��B8/����a������&�&rҪ�|M�.�{������,�GB�/���-��<�Ѫn9���5l� �gff���S-�8tj^�\�|��v�!��i�G��ܐ7a�����p�ef��L)�՗�$E�gϰ�u��mz�� '����SL1I0�M�G՟Ϭ#�����b����G^�$��uQn���fswFj�f`����lƉq\��1�Je�̸�]m�i����8�0�F(t����H�љM��1�5u��IW���#�{�fo�O����p���#��Wl���x�1T7�l{``�Ǵ��Bk��o�tf0�i.��`~  ��>h����6��*r��U}��QXXx:�"�]{�z�q�_��՞k�sa���2�����/����@�� !3�L��p{��f-+���D�Z<�]#��jr�y�驩�2/i�;LL�D;�57�/�m#�h�Sa�KHL�]֑�2w�/�� ����Z\��I�W�7ݰ�hӟ��~�*H���8�OɿA�hP_��k|����g,�N�)U�MI�ە��*ܛ96��/��B��d������%TU���W��uՅ��ST
aď�)aI4p
Y���v�߂��9Q�i�#�+6=�V�:`K�;a!�?׳ޗO��no[Ae����i�	�6����ĝ��&��������M_P�V\���n��yyy��}K����D�}�~�����P��{��^@#h�l&�������;廉�E�pݫ��`׮J-,�]�5'h1�(VI{�2�ూU��#f�3a���S}�Q�tl(mc�f���`MS"�>�~5�e=�@Ks���=����j���KQR�A�uW��4ך�R�n�{�=9$O�|soϋh}Ua�ޏlBe������99������#��4>Y���z�L�������%��)�eE����9�iшl$̒�'mW��|��̡tW���\�2�t��ns{Z^����٥��k���Oũ�{��\�Ə��L�h��r�?3Ĺc�Ԅ%/���`�F��= �4��r�x��t�H#�U�H7B;��̺=ڮY�(�=PM���L��>����Ђ^I���|�ߒ�a�3�A����ڵ@G�W���К��z�E��׵���;:K|��~i���d��E���b��ۭ���*S^}�Z0�������guRRXS'k.cc���8�z}� k�%����v(�ڍ2�d���&��m�e��P�R�vq[3�N��ԋ3�3!��8u5�É�6�4��n� z�}G�a֒��yc1_.nJ�V��C�o"�S���7f;�ӧ�\�5�4L	������A&g�~Ρ��*����Z�ٜ�Zu��+\4��b�Nc�F������ޙ�|�����R�1�3sԤ��1K�1E��+֊�����C�w.΄c,}G�9jJ��(qN�ւ`TUS[�u�i����T������[�#����0:�!(ck[�7��<cy�з�̯��N��qOO�徔��i�գ��K��$,�=	�����ә� �Gߣ�q2h��R�6�HÝ|�/�/�,�a w=���H�A���;m�|�#$K.æQB�����0��"��#�;�Շ�_~��I�h�R�|��̋>�"&Ts���'��̣@�F��\�[��a�[��冕Z����.�8͵��R	���:�6�J����frC8���P�~��Q��ɘӴ׹;L��>�b�s����feϗ袕$�����w�׼��x���Hf���ˉϷMJ%y�"'\�X2�^�B��
���{�Z	6t�A�>c�\�3W{���+r2�GnU�,##��6���f�;/QQYٲ�r^^8�6 �SSF���Z20�e�������}�L����'Q�ݙ���r�:�k���<�������-��~���JK3�ѭ����E^���GL�^���+k�$��i;��a� �Ԋ
8S��1�K~����n�%�+����[��s�-�]���d}�F?����hi����\YW7<4�I5�KLl��o�A3 �%��q_Y�P2K6��h�'Fk�l�{�dl��� &����秈�?l���mL��;�]?��2���4�J�Hܩ��A�cu�p���������I�Eo�+T�s�-���%���\}�cag�1�}$dt;*����V���)|4���˚��2�b��-޸�8$�c�b��<y�o��+��Q���B��F�k�w�m�<��T�O�>u���P��5�#''�����@�ʊ���@��p�Ǧ]�F�9Da0OGIG7�G�]�G�f���bDf���g@������5ϲ��[�4v�&?<	�Y<k��g(�u���MXF3et���W<����%�����>)|����Lã��]g�����T̰��8]�t�T��\�	%e�b�G��V��P�E�M�@ Jn�.a���w.�{�4'yS�AB������W�K�?�ؕ�R]ܾ�x��r���8HF�g����IX���g��W�N
��e^��)Q�lQr�����k��c��CS�6?ڴ���U�+B���E.je.R�M'9���^@�F1��l��`z
!��8�oLL��z8�V�qӆ��^��� ����CJJ�2���UV^�707	���+�������*���G�{����%44ځ1>ٞq�-�?>N���wQ�U��>~oX���Q���c�I��?������喝��I�QjԞ�B�0j�Ǐ`�8����K�t�ӊ�����~f�� �e������qK ����|��|r���?D��O��Th�[��b"ʔԬ���˽���y��L�d�wOr02���eB����3S�L]����Hj��˻:�����Ҍa��%���6�S�5p��X��D��ê�5�K��F욋��B�&��'g�S���J����'T�����{�Ԭ�b�)��o��
B��b{S5�2ql�gi),�Q-,���P��[Mr{������b���+yy>�ԑ��ߑ�W3cE!h������)A���eM�{�C��B�p	�A����^A��w96Y�Ⱦ87�k?�]w#4-*1]]�>�E|�JC���So~���{�^����Z= t��L��<�'���Y��ﴏϿի���(�\J����,�L�U�9������?T�K
)�C^�`M��Ϧ ;J(á����5?�r��yXo�7!d�!**T���%�'�LHv�Z�d�sՇ��Ž���3�C+OB���	4oL�����g����3��uW��̹���?Ny�z>�LO'��M~�.:xN�U�H�M�1�N��'�Z|�s�ovl��o�"�χ��$�%x-i-5#�f�'r�'�$�b��������o�����oGJRDB^��àr!`�SũV�'k��ЙŪ��3����x�4�Z�-X7���({��)�`+�`�Z���N��K��E�K��ǚ��(�*!5�e�D��xQy]m��c���䊖~<j�CG'x/|��E�����˴ՙު��!����G����5��O{����Ѵ
�>��~����%����s�.�����̃_i��jz���l�)Nc>����s_�F�NH �:4����+��P3230<�!`�!�Od(V�*W��oGݶ���(HeKJ����6ڟ�zV��&OJ���0���m��z�-.����g4���ǎ����i+�[ ���H��Қ�|(�Ց��.4V�:>.n>����5 ��H����y��l��	KYGG�0�ƻ�l��>���X|usSآf�QZ��_@@���3���p�Y�Ռ��~=��r����t�Ջpi��W)�a�N��ncsLa�"�p!���uH5�K>��z,��������C���,����M�s�����%�c:U�nB/~x��~_"Ǥ��N��h��+���ȠF���r�~�jH0$+���@q��YW,��{��*�lS�P[�K�g̊��PH�7�[�!������~7Կ��ύOB�,����*�������	4��v�JD��d���~`fF�[�Ck��r��y�$�ֵ:�����S[ɇv?��ao߽�NN���'�hUw�'�'�?;;���G�����F>�}7��hhh i��-[����	5�=�3 �F�6���>�#,,�9	���v�L��A���J�(����1g���F��:a5j��?�����(/��B�&����r!&J�
��y�wNJ<.�k������e�o�������h.U�uJ���wK�8,-8�?������	 W���MM���y��Ӭ�R�ڴ�۷o�'&\��̡ҵ�������CWLL̗zz����k.���Ձ���\	u��Ӄ#�>��M�G�{g}^�I�!������G����Ñ��S�y�z~q� ��ۑ��S��,�%���=_���1���fN]��kw!ܯCƨ޼�|v�F�-��o	���5�v/�_ݵ���V���)�ac�����5{N���a��m����v:�L{J5�Dw2|\ѧ�%�*��Ü��CThT�^ ���`��D1���U�1X�O���^U�|����f�[p�`�qd�P��xx)���T��>zU���K���h|��knβ��b ���\�ؐRT�-x�&Ku���/�ܥ��-���N��7H��I7[�h3����n�j4y6$��� ����`���m��r�ׯ��� ��S+	ߓ'�Ӱ�]'�8�<���@
�@>Q�_�A����G.����jU>Q⸥�ܠ�9^z�G��#�ѽz�
>�S�x �4�;?�������b�w{�n�U1}xN�V����	��a�K�;@�N���72��DB�8��G���d��%[��e�
�T���@�]]Ǧ�y��8 : Βn�����Ӹ`@x��GD�:'��GD@��:�����FFƚ��B{�MW8J�g��>���o0����1�]�_�᥊��c����lM`�N�
���Q����M^�w �O��"'(*++��QQ���M�Z�Գ�$?�=�z?a�I�ug;���I"?��3��r"����#Wh��G	`��y�����t=\���dddP��)^]9�y����_�9ƪyg���?K�m=����?�%�=��E��(_opV�3x��G�ϭW:�C�u<��|=��| ���z*���J>�ɛAH,�{LZ����eT�>[�����w��9�����B�°�y�t�[�4�������6E߂�YV�>r�sJߋfm�h��� �ST����B	���]NE�+�/�-%��^Wb���;0G������̌�R_�i����Xm.���j��ni?)	w;�c�����<G��pa�|N^����yI%%��+�	�,�%S[�VN�Ɛ���=�2r32��yB��Rϝ$T���f����aI�����eH$��j�:>z�]N��Bֶ%-OCغðУ�]��g]D��1}BBN5����}\|<�w�GiلeHJVV<	]��w� ~�VU����;��zs���|���,�<��Qutա��R�K�D���%�j/z��=��W/6�AE�oM�w�	b9 ��O'	)�4b����$��F�j�/�R3R�O��ÖԞ�f��v=w����\�M�uc�8��H��LHϴt4�/Rbo�쬞�DZ��N�O9��_(��$�t����N�5y�Gc+���e�'���҉�ЂBN��$)�p�\���`�x��m]Z,hck�=M*���m�a���3*%O~��1A���t����P,|�Y8��PF[�dYi��-�»�w �K|�g!�+3�A�%g8(D�FqS�8M��Z4������||�Ư怣�R�RTn�� o�5����MM}���X�y_�֟��^�-�H�锁�x?o'ۭU��������߿�Vd ק��ze��� Rκn�����>�U��[aҤ y�/�Qe���Ҩu焎�P��ǹ��L4�ė�'jpF�މ��x�M��q��h��tu�/v��s0w�� N��EP|=��S��SY���C��Q�-��||�E*���j��a��0��Hˍ6K�PIE�RRZ�G
P �972_&��ѡ!��9O�<��3w�$�/6ˡ���O�i"���������d��Lq#�\9��b(s ��+�� 3#���X:��7yrtl:@d*�72��P%>Y�s�c��!�n|�̸����4_#5��4�U�+��=Y��.M�g$�]Ao�4�&��_��0!�ƦC䚢�>.x���>P���9��D����Ϥa�;����ϳ����O=A*Ey�E�6��Q@JrtHߗ����4C®��Xg�W����}�m�w�5̫� /+�7d�0����KE~��_�wL���	 9JO/g?�����sW~
\�7o���[�����cs2��(�$�p~��K�?^.�ZקK%� �� X�2��
��S�z#
�ѓ3�����	��v��GO�M��Ձ���S�˛C�եS
}�97&���J�{5nR���W��W=��hW�bs�Omv.)WR��v��w���A�V����B\\6ߐOV���*���e���>��&h�;�����S�s6�i�вN��L!]S��@hj���'#W�Ѐ�r��q�?6�B�'���RF�ݠ&�e�ѭ���Ӕ���=���U��v�ٍ��qq ����ޡ��&��/���F{=,;�[[%�]V�N/W��R����]��7�g��TS�v��;s�c�TΚ���n��P8`yM^7�8'�������W'sr�h��J�?H�4a��eU��Ed0�(k�ZW0PQ��jDի�*�
s��:��-�9��2��5��}l�f�@�huk+i�I��u|��J��I��xER���T�JI�̎�F	1ƕZ���r�ʴ�ܡĮUi����G ���#i{V���>Fď�_��1�{���m�8]]�Uh���s�֛!&�����:��89���YB�~����x�ص@\��N�		h�NkQʘ����� |����8���OU�`��M���W�k�k��.� ,�U����ee1Y~ol�*��7���6��FKZ�P����բ0֏t��O�g�pT�����(�ƀ��.�	�ĪP+�)E��U<[��9��m��<�k���kg�1�q�vS^I�r-���3��DSP[QsSٞԨ����XF�#��)�y��G���Ma���ש�4����BG����%egg_��	�t����fE���*�C�� k��SS����or.�{�5�|���8���?q095e��Dk���x]�m����*P]]]�[Z~;>KOO���?��	��y�/J�C-��[�1g�󡶝8U�`��e'I�4E��(I��}]�.kЪ����Oq�c���������g���܄�,'|��%���2�3<�}#��a��R_���I�e�n��8]0܊���ö����4�F����!��tK\�0p�c�$���;�6{�VqRRR ��3p+��!��aV����7���x%�ܾ//T�֠��l9����������DI�ﾗ��P�h�D��U~0��	�CiN���>�Ϟ��7R�#�G�q�#(�
-@��6���%�_o�Xw��w#@#�ۭ#�� �&�ߜ��ӧ�8O9e(N\ӫ_l�l�{�I�JL�	
����>B)�{�ȟ%UB�Sttt�L�&x�%�G�w���X����^���Ĥ%���Hg?��V]B�^(�SB�"�u[�P�4(	_&��q��m���y�'�4�|�٨u=K(T���qk1�W�WTW����l�t����*�Y>Q �.�C�UH$##���${�ZXI���n���v xП�g���L�d�����D�r�MοVF����KW����fT:?m�0c%�wCy] �RYYY&*l�R���;�f���#1���̟�]�ޗƱ�h��-�|�{j��x'z�����2|�ݏ��Xh���-d��_�Bxe�(�p��L
8���������;��ܗ��C���fD����k�
4?C�K��Im��`������ ������>-Ï��f��#X��#��#Lp��_[�� �9ӢJ4��� %lQ-�MY����lmm�Y7�%�m[ �CH�P�'����p�\O��7�8��A����=J��vz=v�ڀ��Qn�\M)��';r�$�BY,��Y̴��c/�eM{u=��r*S���/w%�x��?����'�x7hK�n�>�2c:���������a�γ��%�ł{�V���(����GAW;�}��̛��)��?#��g$Q�Q�|n�n1`�~�z�P|ͽ�vR��,�%y���4dd�:�y�}f�D��x�_����ujE������ �ml��s(F3܃�]�H�'�U��Eb������@���ݷ�2<�������2�t���i`��7b��jj6�d �]hb��8?o��uT9�2�7k1���"�$ l��E���4��A�\ �^&���g��_3"���?NA��q�6q.��]R$l�Ψԁf���1�0{v��^��<�صC:���$��E����u$7,�DB*�ŕ�S-
V�)���q���\�*JJJs+����Ϧ5:��%a1�YO��m,S�*c	��8�G
�&'S��_T�����!$�H�L��q���%��	�N�GB����p)���O��̀S�^U�HH����v-j�VvW�w��V�-��N��q�����*���<��O�4�i����ލ���e6">Y���3>����,�_}�6��i=;�7��o���e��t͢'M�qy8�2�Kmq�ts�Q|+���,��o��]��9���������`E	��)S�������A���f8X��&i��w�Xo+Y88 a������2)t�	���iz�z"
h���J�8݋&NB���� �>��Ihkk�XY���s�zG�o�o؞e��n�G���p�$䴸�N0�w�9�<��A��������l�T'��)L	�I�*k�����T�h1�l~���|�E7��ۭ��vE�kb��x���Nݦ-`���(�\Z����ص�Z�"*<͇�J%Q��لݗe߇B��a���Y�>44)B$6��0|\G.�0�R;ne�}i杚.(]���"z��Nf��5]r!�Bۢ�.�:��z u(����5�K��w^y��mU��N6�no{6Q�.�455���	_>��[���N��
U��4ݡ��ݠ���[r?�W�w�HGO�P6��~����X�n2Y��.뗗���T���a�.A�w0�CT��o��ıoQ�����e=�0x�����L��G�P�
Oۖ1�m��� 
:�A��EB� )D��0��ChBƱ���}?鿿o�#����6V��{�i�@0���_cY&� YH�"�������B=r(���;)����/�L�gb�zY7�� ���@�=�(N��D��d	Yل-�能=O��f��DW��_
0�Nǭɀ�m��s�W�,��,/M��ܙ_�B�����JV���1%�d�K����NNN�Bs�)�j�MTFR��ߣy����UWΣ"H�+���=�Mj�W�Qiؕ���|}���)-��ʂWՠ.���^�F��i�]�H�;	�3nkg�� 5b��EH�A�\��V�K?��H۵�H��v�~��q��?R��O��ښO�A��׹�����CUi�8�
�Λ��4����t�tCɛ������r)i���L��H�{�� o�|\q��?���~R��鋤��1������ mP/�H�T"��- G?5.g����q/෬��o � �7�!���%`�?�|�ص ;09�h����0�r�4-ㇶ\�M��IRz���Wl��I�?o�p�k�Cϗ�ME5��K�6��%��}�'??ߦ���ْ��"\�2 ��ޝ��&���t>]�ߦ)b������	���8w�]!*�@��Z�E)Z�equjG��0c>Z��%�C#��O£����B;Һ�3�{P�V�Jr[JU5́o�_�=�����Z��Tl�Eڃ'���*q�"+��pqe�{�F6z��{�Ώ6lk�����=�Q�����k����Vb�MǕ�A��̣e��E��M��2��W�,h�A�Wz���"o��������r����r19�R���
#�#��F�$���)4��vb��wE��1-G��*"*%g;�$Š����¯�Y����MW[:�ܨ�>�Z��9;m׮,f%Z�tq ��0y�:�ˋ}�����y��O��ƉaRT{֋��I��To�o�V/٧9�nF|����;����B�8�����x882	�����v([|Ѡ� c=QĽ��'�CK:���i�9?%�y廯�$�D�7%l��W��l�JH���|��J��8�	��@��x�C�;�<�>l��H�,-�^�k&j�����s0ʷ>���/���9���eb��U�(4�쥈o��a}+m}b����K�0�t��쭈ݐ�"�3�+,�sq���@v)����ާԠ;c�:��d��4H3}�D�Py�K~���ǒ �%j@�FR9�oN���7�F���COA�&�˗���n�~Q���ݘggg�mi��0+�zL4�,I������T�6��ۻ�U�[4�"k�/lY<�^��Yu_����hQX�SS �xr���%���%�D�F�mPJ�-Y}y�e�o�p����)�P<c�	Vub�ٴm{NQ�uA�)�;�-!8�@�8:��p�$��%6�R��A�~�����4a�"�p%�=�KO1�[�_^�ʃ�j�����9̞ˑ�䃽Nj㡬 �B��o����Es��v���,�$�������<|ͨ���r�Ho7>���3�Ϧ_z�st���ix�����Bs~q�	�S����5q+���3I�?��.��N�8�F#��Y>�v�.���ܗ�Ӣ�/��R�����1�E��Z �'�
�{T%���_���g� �U��w^��` � A�-Qd���1��/^VV6�L�TE�>��!��Nyp����c~~����;�>}z�*/-�sbf�S��$#�f/c����h�#��y׀�5�d	dt���7�����"���!X����.W�m�M�,�:�S�tg�z{:eȒa�{�=�^�v���2��Jwm��0�����X}�BA4��b"�F!�-�İx�
͇Vڳ��h$7X�Z�H��$����	
_�n)А��iEii�������fO>�����A�2B���kH�22 ж���8!��2�^(/�����5؈��<���r��z�\!&�]����<�*N�@5L5���[ �}�,�o�p�ma�p�糿�mDy/2���!�4����h'��k�����M��Ԧ�����!cQ�L���O|�$F;�1��"��Ux�Ɩv�B�c�@!�ЁZ����q���CY����s�Y�Cj9���Él:(�O��ѾM��e��&�������#���#��b���_���E�^��i_A)���.R�o��eNi�Pt�G<�aۖ��&+�XX���������^3) �L4_�)�)���#yj����!PDh؜�y!����>����Iv�R�Y���������g7w}Ij���[�=j�K�$%%e�E0�,�f=��:���񢍇"���w�Q��X}iXj�oj��NXL7� ;��X�p��f��k��7=���]�v(>��Y�Z���%������G��߭���Sp"	���ug5,�W��?m5�h�;C]d���<���ք4����|j~�^�5
<�qV
@�p�\#jIn�#/�o�H�cf0ڛC2��� Z�ߓ�	����U0���_�G�y��O��|��;�'nН�� ���6#bB�2�>�3���X>fw�]1tGV�)阮�h�f��Lh7W�vN���J������7�bUU����PQ������3����]�¯�=����ɩ�iN�����ᖌ_=w��ώz�"x�s�|H�VK���,>lły[�:>>��y4�����@�Aw��2��*�4��Iw��<̂��]=�,�9��{	�Y�w��{F.ݟ�4����`2qz�8���03������ʶ$X�b	z��:9R�_z@0�:!���������J��ŉ�j(	뺩�R̝s�C	|e)�h�~��pR(��İO�|���Y[[�΅��{�	��4�`t�����*�(�AU#*�K�n��������@����%��uP�|6�.��pVm)�ՠ��t�(x���h�\O3IĐ�e(9��C�L�ٳ����zL4��7��2I�l]E�嘛������y�|�.��\��A`�;�'g?n�����&�_����I�S$�̘������H�?j>��ʧ��HJJ2\=�g�a
Y搈��ʍ�MmS^7�J�����\���1o�"a�#y}�_�	2�_6�/#����E�[�?�.� V�����[I��`	eaa�p����ϛ����m�[�y�!��x|Z� 5���9[�X��:�,�?���3٠)��u�N�Z��\�T����2b A�����#���O���",�ۯ}�"�囤ǈY�jϏa�-�����͑<BQ�+m��O�	����9�#��2��Z���Ge��RC��Ň��O�	a��P�hG����vM''>��5GU�@��4�=qorZ�}������F�Gng��9N(��x������^���ǭIJ`��g�T1���[x ��t�R]8�"^<���n����w��Z����32���
���,|}�U�99BoǠ�.Cu_�kA#�IU�����qG,u����Wz�j�>&���*n�>?��s?�'3NK�^�K�R�tlӻ@��GH.=Е�I�&e�*-K��vz�=$�W�LO�M��WWb�y���b�-�)̈�B�=//Z?������I�m�$��` xi�P�oKvdm��t���	��qFH8�Uhݑ^и�Q��>����-��L%2�ĳp��´��N��]׆��⠹���b9�N���/��W;^�"n��I�Q�"BD��5�@'u^�* E�c^��ί&�É����h�z4l��m"��B����x��\JA�5�78XV�Vs���!�(�� $]j�NN:}Z%N������#�@�)'�����K+��|ݙ�����$x����������H�͜�}��oi����i�>�>R�����1���z?�(�>}Z��"�]]��뭭[D��L����@N���`��;�(������y�Ɔ�\+��.��2/v�T��BѤ�zT�O���fW�ݬ9fㄵ��v���0�D��3����qd�<P�o�݂U���L(�ʔ��*c�Ujg�z���v>$3�}30>��<4��O|Τ��9G�{DUU�`k�� �U|����p]]]åc��qi�n?ړ�8�[��qk�g$7��(��o��j1���>E\�ɿ	w����F2j�4�����m��3�
|�ۀ��"$��UҜ�|�HN�G;1��]�Md�����r냗��quS�������A�����?�z�/�W��5f@�ˁt'�x���t��"�0^�Ǳ&LGGG��ot�9������gr0�5�5;${�!�t9�˰)�&9�0�\%a42?»�w[;.no�D���ɹ�@GX�����ι�vk@��B��F5'08�ő�V����u�۲� ���B���PVx�[JY�?�s��'Wb�1�S�y'�e:96��ը��Ą��fƬ<��Y+��(&1t���]���CE���v���C�U(����ȝ跸o\��7�\����-/]�m��F����,�e���r�hp�Q�Д���;�e���}QN^?��5�@8�L�@gNȱ�}���l��eu+�2ʰ���{��.������n8 ��88-+��I���Όv�l�+9Е�ʖ��$��<� �d��0�$ۖ��c�S������h�[�y�H�vY9�S@�����N����k)�u011�fB��7�}�n���-b�zq@�z�d�k�~�^X�߆��{���3���H������%Y��]��F��[�K���fq�������%�KP2���E\����e1�f|+�E��Z���j���P��-�ׅ�������hDD(�I�1��@��a�3Zl�K����hd��-}F��'>���"f��(2j#�L�&�50�������œ�_�GHGY.�C~��}_���h�8,�+���N����^�#��P�YZ#��,�д�R�3�v�X{�N�q�?��:����^RS
�;r%����o��wN������h�M����7��_;ȗq�^��j�V����mya�`a���!C����Vj&@�fJ��\\\�O�˦�Cc� ��-��{vo�+��~w*�K9 ��v�۟��(�W���%��.�O%�dY����50@��C��E&�qq&!�A��=��gԮ�y[�8��AFQ�]�����	U�����60m�k(|4�b�G�����A�A<��r�X�/�j^�1��IH'^�C�O�z?c�,c�^"��cMF��,�j��)lQ��z?@�b|s}�a�͎T�� �m�)g8Lb�,���n��:vr�(�}�{����ô�,��G�"\\\�	O��
������L[��'� yi�K�A��@�?���6g�%b�x
��vw�m��\�㋧��bL���ݾ����8���0�	�ݽ�t�賷�3K���-88�#PeKFCC���A�Y��k���r5`sW2r��!%%�Z�����3u�Z�D|��w01[�^���}���v�NU��s�g��x�#T�;=��x��Atuue��58:�I�]=�H.
�-�W�E5u1�Kn�S�d����I���}���9���k���[�P�ޤ��>��t���ߕ���⿚���gb/v]�a��b��yh1`P�Y�^ ��T��ⶈ�-����ϊ�K��oZ�=�aZ��L��^V�e�Dz�/..ʷm	 ��j��m+�J�.Z���]_��+ t���Zz�|��ML^�y�|os�3�����,w��승��e���o���z�#����E�b|Ǆ�������Q�XG�`�7f��Wh�ubY���	X�3�4��;�O���g��pH5و�-�r�b�`����Ս��vR����>H����N�A8}_�aT�L>�'��SS�]Q��a����)�!4�VY!����y���!���ܴaY���]��Nn]]�ZF�fЗ,������7�]>Q`�	�<D�+;}~�İ�P(���N%y�5 �n'�@����d��})�x�]7
kNf�J?�5�^׾�~�Gמ�����9�x�S��T��o�]�l���d|w�^�$��*|&fy��tϞvQ~��1�PQm�ߣ^E�t��tHK��tw��t34("�)0�t� -94�1H����^���b����y�{�s�y}2�Z�ms�^0w4AHL�QUE���՚Wwl���P^^~�H-�r	�:D�R�@��|%N��� *�C���mS�����A�� ,�w��c2m�g�����N7o������ò���,�X����- �km8�y]�k�������gO�hi�#`[\���"b�7h럳y퍾��黗����-���+]]�]��m��M���{�j�����C�}+[��SY�Ι��Ϝ���?Zc,�y{X���޾x�S�Ë
�h�9U�n]��A�>�DVYYh�,��:w��=%���߿�G�0�@rlb��Ϳ�����5 gNc���������B�s�{{���(Y�����C1���!�9�A ��ɉK����^�5�Jo��#SS͓�o�i����P�1sy/+/���!bz�k�؊�/ݽ�}���+�Fl��:Ek@*���� J�}�*��$�mU��K{'��cQ�֢���P���.���&�i_�� �_g�4S
�X����8�����p�{6�^D�N�1<,,������T9�o�z��r����(����<���$���RUK�ᡡw��$��`C�J3�)��cJ�	H	ş6������f���'�H+���ΐ^^��rnT9�����".>����uyhwy#��5�'�[������E����_[X|���{�Uo�����b<��%�ՙ��O����:�i?>^�M3eѭ�!b}�P¾����nn�Y��L{���"�GR��4.�M���⟒�ƽ�IL7�n�EQ6,��UD���Zj��t���-����6==�ck���{P�۾��9Q;nF�	�l�k�P�qXO�N����TM�>0�:��Qu��!�����E�L�-����V�2���/�k>,�3�$�H�Y�����~���5/��ޞzn�{^<*����K���č�T_��s���b��5vx&hY�>B�t�+.�|q�V��M�vf����;�/�У�*�f¶&+iXYoC�\�����W�`�>�>�j�ƠH����L�i[]Rj�`�h��/Dd�G���'{�!���jñk�^�ץ�ͪ����;MF�.���i�RDf[*��(1�9�y��5)YY�������w�c�0G���`�۪�JRű�4�di_�t�	�c�&�֍���ަϦ_�2���X-c�ڵ��B�[�����}H��?0?"d#{���<��t���5�l��e:Il+�X��bt?��ܨ���^��Ds�L������)^W�c�_'���w���ձ�����m���J�û�%[:����+��'��̳���c�j�O}}E+lQ
t+��8��{��ʐJ��q�څ"�3��Уe/0gs{=���Vo�AbzM���'�A�7�����a^އ��R5ؠ�c��+���}��Y܅@�Ԕ^YEŋ�gK��!	�A ����nQ�n�xi|��8FT��F�_7	��L8��c��J��/x�}�d6�]&q�ٿU�|�u��U�@��b�M��BBcbbn���`����ҧgV8�(|�{��_�������>�.��Շ�����GBz{��j*O��F/�]�	�����������wo���ߡ�ލ��`O�DebbY
����*ъ������{s@��u�w�+�����;�僟��?Re���	^�q�q�|����e]���|��[���~,��IE��0���E�]S,���=22%MM���S�8�L[s[Ҋ�_(����.�����J���I����l��O�b�AmI()%TU�ǣX�@{ʐB�~�����z,229�7�u(��~�0(�le~&2侥p��!���5�k*/�$+�o*"?"���]!�	���WRQy�������@����?�L������z P��*r�Yŝ���T`0��m���bq�����̎�:���~q1�@+3�5������'�i���@�*')D�Bw����
J���n�m�����-�Px�py|�X�\d�;]!�$x���'C?�����b�p��5f2�D�b"�#�tX��]����e|�b�����pZ�f�(���T������0���3L�g�]�����a����ar�����Y�x�3Ӣ��ܰ�_O���qG��mZZ���p2�cE��U�U���Ó�r���	C_x�P�=RH��&6�R~��i�Y�:��ۯ�A$��~�9P,)H����L��k���]I��^��'5�	=�������X D6�x��s�Ҟ%��D:�ë)B��$$$�/T��-F��#�L�4R�!����Ѽ�������|5�)��}����1S�K��h>�/��H�����:d|��f�b>83�x�����̬��F:4��� ��P��Ʀ�� ���۫пTWk�џ��"��!2��t{�Q��J�b����?�9=�j��p�-��6KO�b��):�[��>z����N�	�Q���)?^1ʔ���XGd�KRWQy(�)���g�a`�ê�EnW��(r��*}F2)�`f1U0�4 �Px�i��[6�3m/��K��� t?�>Ya��E|��qq`�MMLXY�)���
��o���J�_�;iJR��ϋ��@h뛛jpxeMm���t!��iQ]]]uC�"��Ng��?8�rf�7�����unO�zɮ�WM�2��=��^"�N!�bd�|����k5��d�<�
I�6�IG��R�?��{�}]_��;Z���c5.V�
X�(D�����?��σ��l):�2�&T=ڪ� B��:!͈��щ�i�f���ɂ�\&W��^����{�]K��t0#��/2N��}�V�L||��r_��əut��
>S��n�1R@Df��%�0hV�1�?π���P�vS`����I�����3�Dyee��W�u3�܏|��f��[��Z�܀ݻۡЩ�D��z��icfb�Ty��q��9?~)�ٽq`���P��uī�_�|7�lϫ���q륳Z�9)���ۈP��3���o%m���h�iqj3R��Άݵ ���� |�����$+@��g8�Q���U�\����c��Qwy���Ht�{}�6H����=�Тmt��n{ز�P(�.�����	����\Κ/x�W����}��|���S�U/w�,��n5�Â�<2g�RI�w� ��ڢ��Q�����,����S���8��Xuʠ^�u�R16� �P�3o=Q��=rM;y�����%�s�s^h���h۞bim��\i��.;XP9�+B����%$$�^�����R�F�����bx������Q�� ��>����Us7��g�=���Ū�k
�D�����1.�'�Jj�SO�����y%�tU2j�;t9�t1FT��y��,���50��
Li�_����*�N�\dOT�V�U����Qt,7�7_d�󩇷����̶:;ܒ^�_��355�̼��������Q�����z�B"�����`xw�j�����8����쬈>E���.A�5����-:::��_��M�lUL���L��dq���	� �4u����N���>��� ��,��2 �QN}§E���!�Wa0�w$ab���V��=��L3����պ(��!}O�t2��|�B�z/�K�C�L����e�a�R��>-��3vm��Ѿ2{e���nO.��SR�r��!O�A�����bG�KQ>��2�x^�x<j���p&�,�n|�%v��5��~������1�7`�[0V0�d��?���������p�ә�m_g��$���A��q}�O�!��JJ�G=�{���F��0�tv�|u����E�g�k=|3e�t0�{��ޏ��N��x��/j��'�t0��'����EF��2>�%�3"���,�����$,�FX�7���JlW�����C��kF&iPV���ѽ��ֺ��Tac�}}o倴('G�ǧ!��i���#  ���V�o)�>�.�8N	 ��v)^")��8��ibAC@��	�E�;�a��O����q.��v�Aäʒe�sJ�d	���%���\�?�����8xr�.�]������B�3��p��j��{��-(Pם����ܗ��8X�L�m���C����Fn�֎�f\]�Eտ�Ю�����D�7�:�(�v=v�d�F~uS�~�_�A���#��uk��1M��L�n�:����u��c���[���܁$=
��;/[�c�n���a9Zk�iu>?v���yd�B�f[��4r�����OH(Z�Z�0s����w-/m�K��T��fi��g��B���k-��j����� 3���h=�VB�w�d$�П��/'^�M�IMY�ܛ����A ���y��+w`�!������1��|v^�l-��X�|ζN��Rٽ�d?��[���8"ǧ���<cI�O.�8hZʾ�O�����������8�S�?q2KI��x����fPV]C#(�������8�㜳+����t�e�v��K3J
���̽�~��4���4�IP����*I,�<��~�t5з�BT6�����=���@���V����Z��ޓ�1�ꇋ|�y_��j\��#���a��È~`"+l���$--=�{�ʽޠ@��y1����g�pD����?Ж�vSqʙ�V"�����>[B3*Η[Z�ǳĞ�0_."�ˏZ��HCӲN�Ҽ�@<��B�B�eD06:��lZ&��Hx�ǽ��
.3���aԢ�	�5� U��!1fă=��AR��E�S'�d�`j�����F���{p�����~��f��s��M��mo�m }�f_�߳ �Zk*/J�b�ު����?گ��[�S�����dt�K��r<��5�`�&IRRr�jtC��˴�N�Ѿ��~����v���~�}U�E䨺�s�H�xS�a��T�ZU^�
_x)tӻ��|T%éԹ��'U����+5q�$0�}o�b8W���E����x�S6$B=CV���L^�-��خt�:��\\\������+�i�2�HB���zD5�� ���֮��8c����%A�B�b��T"׈�q��UQh�c3ei�ങ�.0��r344�^w&����u���[-C?j�I�,���h����l�4�?�SQ_m^�K2Q�:�=����{��e�qT���,�_�S��l�:_��V�����(+ۺ>L�r#��b��(7W���jp���9�Cv�(zőhM8���!x7�M��`c��(� �[cq"��	�����[9p�/�R4A�Z��>�`cc/��`��%áU���Rpd�<��@��t�ϟr!� �¾]��槑|��5R����|�Y��3"�e[i����"r�yTJJ�z�������N���B`0�us,����g!��Mj��u<����̬����ю���d��OK+��AY���qk��`z�A\�W�9{N�����ard�i-��Vt8��n�N� {�xgAZ_PXX�˼7�s5:""M��^�v�s��KT�!.��s��}Qh=m����Eej	��-�2h��*�����:�ؕ� ��։Rs��-�,Mw	`�5�����F�b��9ԫ,y��Q��^}L��ᑑ��%.NNn�Sg���!��k���3u@5����K��4�󊺎�/,�̚b��QZ���^��;��D���oř'��Z�JUSU� s��ꏃ{M����A�ĕLp��5�M \�£Pb!�]?#���:�I�B6dע�5�l+A�������N�=#,¼��A?�U66�1�k����ׯ^����4F�t�0s�U�k�Si�TgPtq�w95��R%�*7�K��`�r�|m��`�o�*�Ǻ��4�@�� ��L��2�ܧ�a���B�Z�v"�S?Dϒ�T����_q���ZT�y�È��yy��3w����'�z0:�wO
�ԥhͲ�A��4ӟp��;���*]�׳PY��ny3j �A�DR=����2���b�V�ά�<M�e{zz�Q�"�� �.�=��	e���������y���DII	��e������xl��:�.vN�ݡ֐�9�T�Z�����r�=��ֻ,�_�f[=F[?������\K!v@d���A�/6ӝ2���,�N��H�wF����q0��Œ7C�ڴ��_P��=+�#B� ��u��Om+'A>���<v;金H�����>��|NN���p������D��X�O�<���◵>�g�P�{��Keoܓ,������ �����2�����gĒ�D�r=�y���t��f�[�ow�u �c(Һ࠮�~�u���y�=���hy٬�x>�>ܸ���Xj^Q���7R��R�(�{�vD�I���nQZL�X[1D�9�6���CJQQS[�T_�#xY�j��U�*��ط�MI8���vf�e���A�w�T���55:R�&��<�S�!��l��p^U�^ I���;B��{֠��]�'
�|��-�rt��"c��(�����I%���YY�No0/�Zit�1D!��zL~_�����[SuY\��~��o�㿠�y~�r[]_]URUU�v{����jXd�-J ����3d���üx�vi���ޏ��x/�^���Cft��}(d�����~3;�������ؖkO��'O��dD����K��9.Ɍo����᮹o�텹����&rY�=�]�5�R1��/	5]�ښ(/�����ߤ�;�tut|� �����؜��}FϪJKU=7(�Si�x �@2���C/�rS�}�vUs>\����ƕ,E
y���5�6�wȜ)����&�Y@h�yX�`.�D5�jj�����K��u�z�$����N�}���s� �0�M?wbbbz4Y9T���p�ָ5Yy4~�������Z9����65��VM��M��ܗ��l��SDX��+6��Z_=�/��ս$#��4k�^� vP����Q0�@iD��n��k�QT��H��ά��fo</��9��Kr;jٕ��v�Sm��A�4\�=�$4
c܄66�78���^���;[�~�J����\+1��2:g�ZE�l�,�� b�~ v��q�W��\Ӑ��&�O���2�'���5�F��Exb��E�Dk^�D{/7�}R8��i�ˬ�+���G�r_J����|�
��_C���G�h��(���Uy���K�%=W���A���P�[��:	��rtttL���6";n�p��5=���-��x������Q�=EB΄�5�c�2�,\`h���V|�D
��`�[񌞤d��C�I�@���@B��:n'J�	�*~��7'#ø�x��p�]mCԟ���>ꋤ(§� ���<���} {be �K�,����ͥ��O��.K.. ɏ?�$����B�x��v��})�{UZf�=����F__��):ķoJPw�nȯՐ$u�_��}��^�.Lx����#jY���U� Q�w[KA!L�*< Hs�����\}��V�h�H���3 ��%G�DH�7٧7Q�4�)3 #NI�K�FU�^	  h�nk{P�� �K�U��SPg��TPh*��g������٦5F��q4��+)��X��+>�H�prR��yfhiiY��t;0J/^����6b�j3��H���[c�'�T�Sa�ڌ�n����F2,SY;�՛�������c��G�EbAx�������E��G�	�����n�k�R�ɶ���]���;����%�W�-�ٽk� �rۿ�CFc_l)�N�c�����VJ ��|���<�8��x��X rCc��0˂IXUr���x��]�;rM}m%%�<�����i���� ��F p������Gp�4�q�����qk^��FQ4�`�9��c�t����eW�)��\���4�=��������^;��-J2��:{{G$��3�8-k�,N#��>G���.��Q�;BiM�����+Ip&��}4�5I 0,
�a�ĵ�mw�j�N�ҵVb�! �S잩���7�[��-����-d1Y��Æ�wRt�
}��D����C�QZ����~7��%��z��u�GR�j=07�zB��i�	���	��6�@{�S0�+������S
�gׁ���t�+��� ��z�����݄�ֆzѠ��j!t ��J�a/���VZ�L��o`�7�8���y�v���[A&>q�6�����v���٣3�CkDg���N&"2���aecA�d8��^�S�ˌٷ�����-�@|��0T{������`W2
t+m������j� Z����${o#��}��ؗ�YH��#G���������K����(�S̷�v�Y_2k㌝EL�#��K�z�O��#_���q��s3"���=��Q%$$��K�[+#rbl�v!���?Œ�Z��� cRR�z�R_��XbN�\�쬬TMM���h��R~C�*�'�����#�T���wD/r�C;���-�$C���LC#����T'WAWn��/u7hե�%::���켭�.�#M������Z�����Ɨ�>==>�8<t������5��,���-u�hE���M�iM���_��c^� 1��UK��v���9iii3^ �+�fD�b��u���F߯�X:�O�)����		y ����"��[!��}ް�4m{�ڤ�+��եK똾���o�n}o��p�f�rFH@���AZ 8 ��0�����WN9���6l�w�^G�e����o\��5�I�9>�S��8L�j�(��%#'g��Ǒҗ��K�s[D�7�h4O:���|+��|�Mӓ�n�R0M �V����7:�S��}�i$F�ݻ�����hsH�RO�7j�)HN���NJѴrf���
�tI��VE'�K���:�[{%�*�6	�@�#��\����tx�v����ABX�+ /� �Xn�������W��MWw7y��́���K����S�:U�i>|�2��q�vY��d �	J�١�8Q{�cg��<�^�w�`
vP"\,�\[8>���90��rn�j5��?�B�A�5'�	��VOy6쳽A�t)��K��Hŵ���ƍk�ӌ��,���?�� �G���$u���|���		�	=f.��9�U���dCkKk�lfaaaF+pi�f��O�nYO�XK)3�K~�����X��`�]�
�ݿ������N���)��vϫ��L �y�K�T�f �f1RVMI�������۫����Ѫ�/�$Z���ā�j�ۓ���(6���QI�~�۲��)l5�BHDԵ�Ki�8���q:5�2!��
�9Fn}�������Oe���{�򤴷����oa�0�M���4HĻ�D�,��J�EdgK��Q"o�M�@�6ۺ���q���=$��~�PLK����n<.F�"7��~=�5V,rF5@,0�e��茢g&�F i�%�h}h�`¯���$�L$����i���O�����g��q�pV��FY�������F�G��'l>�s��	d�ff���7a���� ������6b\�/��:) ����A�.窥ބtt��-~̒�Jl.ϖ��jq���p�)aI��ǔBnJ�L���(�]Qu���76]Ӑ�����n����0�1��5�8Ӧ�Y`��D������ţ3S����'x=_�A��BTԿ���:bV%ElF]�s#�j�5z��Hi���ϯ+��0^tI��Q		V6��2j���>�r`����m5��t*�A|?���<W�㓬Ivs�b��p�����]��)vrV2�<��u>����9����,yU��3��j�oo7M�P��
 ���5����tx�� 
�ܽ���Y���8�yu����W IݡFsQ�Yڷ^��,���3�����(d^ƕ���L�s d}s�3-��9{�Dl�'&H��!A� KOn[�:�<���2z�`D�y!G�.�ͧ�M���P�'<Y�W���Yz��ḣ"O�2�Q6@���*�,���j�m5
}e�a��􁜇R�3��Zvw��d[[5v���8n��&(*�i�ϗ��>����-(����=�Ȯ=��?+ʝ)�z��/�U�.���O0>�����������@���: 2�9dѣ�s���������>�h��s�Ky�+/&>�����}~|V��{.�Є���S��u-:�S��]7!IRe�p �>R�X�3'}�%<�m\�9���H*#UV�o+�����Ԣ
+*x����p��}/={� ;��A�\ �>��F�2�H�����/�?��׊"�I"i��R_Hb�7�'�ܻ�ڝ�p�#4J����N�cWggg�	{����e���������"Fۿ�aMW]k��F򕽽���AM^���a�{�R:�Ž�	b�Dh�IIyϊ4؅Od����X�qa��
�˃1�!Jx�����D�iP�*�"�C_��*oMU���ʦ��7�����S�!��r��$�@�A��U-����Tp}0�OcS+j��ؾ��K�����-��b�o��I�"{�}�f�;��4�H�:�ѭ���*q�G�H�9�(�8;g�?�������u+��A�o�aݟ��[�W|XF���_K�t>S�$�Q]kC��j�<�l0��~ ��;�Jߣ�T�o-�;C����� ���M&|^�����3E�!_L_����Ȭ��޵��3����� �	�F%���{�Û�t�q!���3c���*������TZ:��br>0��*$���'�5Y���~���B�$�YY��P`3i�^vE�Idu[�D��#5r��k٩bX��x艉�Wآr��c���xЫ��	 q�+��WZ�Կ m�Qy>�j���y$�&�c����i�����cia���ނ�����GAZh�=���_c��ۍ�Е��7�/Z�:�D�yc���I���E5�bW���Q����	=s5"Y�D������JVV��.�� .�0F��,��Lq� ����Q�B�F�"0�����S����7Pl�b-9`$u����^7O�uM​|��6.d�!�֮ϡ�&{!3�[*}y����N���5w.`��2i����d� ��3�Ʉ���lR�[o��H�h���0ųw�{�	B��_P "Ƅ�,%�`�,�<J���S��4P4��xI(��7��M8���:зu�2E���_�Շ%��B9�#E�#H~�k�d}��m3^"�N��"�7���v����cK���)��hI�0���u'���y�eHT�<�k�����s�@�3H;֢���JD��6X�9P�1��������Yr���T�!�ا��HP��0pX���^fg���D�o�&x���}�!�0���n:��Nni)W�4������S�w�9���2TVN۾\�>=ASU۝��$x���&(0M�4��my�8~��,��	O�(=}��8�/�5��`�����T���dh{8�#P)�.�Ϟ�>�b�60[��9%}�7^ة���f�wk�^t���o�ɭ����_xm&2�@ ���YH���T�u_*k3�c6{�"� N��9�ū�/��)L�yX]Q^��/H����)J�Q�m��d�l$4���B�o�0�����v@��X���Tl\⟝<b�|�:X� XvᛂTǡG��9�/���>J��N2QY;c��ۇF��r��մ�)H�����t���0t���Z�hYG�2�&$+���M��
�Š̑���,�zyX0�W@蔘@��
��К�j��A� � W@z�["�Z�T��ߣ=�q����{�	ч�{���{���4�7Q%*�b�IxA4�"�FF4�s�iiϊ�����rsk�}��zUL�s�IWYjV}�����$��vǰF��)��g�(�-��_��i�	-AC
�p�z�=���S�s�0ڜ�
CT�Eʞ��ѳ�8>�m�g>,!
w�X�+�ĺ,�R(H�T���K��L\\Q���U��+߾}�%1�i0f���j)�O�b/��.^vX "z��z�G��ƛ�l����ut&,����FN���@�Y_ޏK��,��KnII�Gc,�J�'U]����x����<A�x��e�篫�\��-M`���e*��D"��F@g�tttLH������`G~�y�F��L�'���^s,�������"cZ�e�ju���U%]��{��`���������:���x�h=Jg���i<I$�r�mmmh�٪�O�4گ��� ��8)ѪhI��7��Ocמ��ר5�O��uY{I�d���Sީ:Fҋ}!�EEM@o�5�9�  Y�i���J>K���S Yy�i]}��03E���^!r09�}��*\-�y-��q##�.E�F�MI���J���~�F���L6��^�aܔS�-/c?�}+�����y~���2a�qE�;�#�FU�Ⱥ��^!���?�M��F��`x]*#��K�A+9R��B�U�ooeA��\<S@%i�����.>+��h��k��Dԧ՟S�QK?{T3��2�X;g�HN��\<��^W�JSV'T�_���p��,���摁�B�!�ȏ����5�.>���qlM����#��n�_*�xSQ��p���d��W��-7Y4���~�� <Qa� m9R�xi�ie5QB=����=�t��qEQ�
�<�B o7nn�i+=�p�ǣ��{��%`U��,��ɩ�������z����99��q�̼{�i`�&�x,��%Pa9 ������)p���u��n-��w�f��Wp��o/�}� �V�,��Q!�������-RWI����q߰��p�F�%�|i�-�9����8<��o�|[q��Ϣ���*Tߓc
�}�ػjN�P)���E1̔��F���]9�E&�����O�������sO;�8��V,.�Ɵt1l��3:�K3�R����ɖۡ�7W|DAa�OV�1u��x�E_�(���f����Z�^��,��8/~
�؊�X���9�Ġ����& $�F��vAF5<ϴ������_��'_5�WiF��>l�f�R�
t���I�V��F	/ԇ!PK���E�)���^�0�����a�xL׊�[�����t۪A��[�#!~�
k*��v�������g�
����������q<Y���-t�4y�cqU����QjT���F�<���d-Z�=�Vn<�x^.��<�۷�G7���(N�q������W`^������������*�Y����Mӎnvb��K�n��\��p]&'���}�<6�w��~��b6����[��С\�)�zQr=^��i���u�)����ٓ{/[���sF�	�4��q�D�a�g�����B��h�Bo�[�����tOQM�7x�k\��?ȷ�T�r�/S�Mci���D/��O��,���TF�O��%�E=ă�h�6L���d1Ԝ����_rl�?%�G�P1�����0���|Ի.!�/���T߽���NE��rnx�L�ѓwm�*�o���G>ky��)��GK��Ѿ+��|��|h����p�BLJ���e ���b�xH~ԗT4ި�����C�a�����щ7�MD\�����Ş�3���'m��%@�dw��
�~4?;rܮ�F�R�kʊ���4��O<]�Ϲ4e�47��k+��3�{◷T�I�%�]��N Z`�Ģ��;�\�ܝ�����_'勐b�f ��Ζ���B�P�������5*2nM����Z��Ջ'�-[d�5�q�w,�w9��]5�������-�O��IU�kuH3�C�����\$9�v��t�>��oJYHL�l�"b7�N6m��G"��>�[۱ިK�w���I�,2ol�E�#���.�L�,��Z�P��&�r~�^4����T꩹O�~9E�v����hQF4	㌛�d�^����������*��Խ<[sԈ�M��n�4)c�..��{�L���h��0q�����P\+���QDQ�&��x�5�.���Y-h�� ;�m}��f5hǄŰA���R�_FV6�F����-�@������|h+h�8\���=J�q���"[b��wu�>+(�y�`jS~7������2Ʈ�b}���@iT;��ڎI���@������8�@��!?��E�lc-�����v�+�� �G��u����3����*�rrh5��Q��b�G�{FK�F ��5�=�^.4�5��v���x��p�?��يHyݷ5
���!���-i��J�Y�ᮺ�	.�X����;m�<kv��:]���`X>�i~���Fo�%���9�7����{Im�f1����پџq{�6��|��tG��X���>���e�p�w�Wm��4+�QA��F<�I��黼�u�lY#|��2�\�s4�B����CR����8�󵊟D���'���@oprr��l�������Q�F�i��uB�\��w+�S�^7+�4+T�~�UT�n-����m���zd���	�MK��*����kI���_�9;ʫK��	N�?qZJ8s�S(,���'XK\�Er�7��4p���~�ν�0����Q=��C���p����O�B���������	��l�������$Һ?�κ߳�=�dX:X?��fo��Ϫp�M'����΅Rqm?���Tg�s̟��䚴�ғ'�����3��FE�fq#O�U9�ߓfii���2�m����ѿ��t�	���#����H��߹nOD3kZ��&�4x=�������7�m��:ar�O��	��Jzq�V��.�����+�V�T���*TO.Umu'��x�k�NDZ舠auP)VfV޴�����b�tW��Ek� �m�g.��ae���B�<���;���ThƸ�:�m��K��2��~[g.k^R� ����n�̅���i�{�[�b����5kSD&qU�X]���-�X~����QY�yk���v��X�ڔXM?jŤ+�(&��L|l���.�_:yF%���f/u��ed�����i[�7`�s�$�91��}�B����Y���bA��d�4��(Ң4?��UHd��q��!=�u[��9����.AZ�i�.�
:Z��H*"kwqA �$s������<�@��%�hϹ�Ȟǖ8X�р��������tSh}�X'�1���\LVz��q/f�*������f.��v��.6�o���(ۺ|�� *6�>wZ֦�D<<�������<����"������M����b_B�(�ͽy�#A@+�����6F@$߾)����1���!L$�(q$(d�"�PV�6��h�(o�(m5Dn��p+���񝳥��n;gf��ُ�V|�GgKGg�11YO��o�ao�Zd�!%�����0���U��������ޜ��wbI�yH\�������n��dVi��>�X螃�GMJC�G]��q���s.&����b~p���@s��@M]��z�GaV}d�Y�\x���$o#��r����".kw[+o��"wX:�pW�j�L�$� �sO}�y~��օ v�=<H�`�Z�����	�\���w�j=�;�0؍R�Q6��FA8zh�5�`HU�e�m��ܪ�L��aQ:Y���ҎKr�2��ۑ�T�d�8�L#��nA���Z=����݊h�������Pf|���N(M�i�F�Wi]�g}q��Ӥ�'rΫ���Ӣ����[���C�Q����(��Nu(�|�D�$��w���S��6"���{#�fa��G�9��E� �tv�:{�H&���'��G���Q3�։���H5���Ԩ;�!m3���k��}�j{cᄅY���?<=�WٷU���5$� �m�KJ`z�=`*̸)Y����Ma����?F���G��XT
"9p�C���$�]� ٰ�ϟpb�S��%
'��7��	�_}%��'l�^^Ssk������A�xu����^;��S��'p��z��z#�W�qB���
<)uR�tø�JQ4�cwa�ɖ8m::�]�r�H��f�F�H����;��D��^��)�t&��ݲk�z.8�%�]����ؼ��~���rK��B$m�	Nf��=�)�ō��ڢ�U�~���9��G�?�h�Qn7��+٘�!֩��!fS�@�<�>���>t�&`~o�34=m���4�V� V7���Ą%�E�ʫw���fc��f�T�0*e��P��5��[��8-��"}�]�B�rt����l6 ��5�gd	�G�q_p
����=��y����(�ء�J�5>�]n��g1pc����z�<Z��i߶�Yf�F��9�.��g�Mn+�HuP������Q��~��_3�;���@F7嘑B�3��Y+'YGfv��~]��n�W�{\.lsy�y���+޴��%��)M�F;Ĝj�r3�(w�<�1�^)��w��M���k�W��}F%my�fc.�7It%�����<��3{�zz�k��Kx�ޓ�C�A��V#,�)�	�Q��Y�;��A@���J�k����EM�ՎX�r�ϒwcԘ�-�Z�@�O�zN}}���
�Fy8�ܝp<)�qqz�W)�Rʄ'��941�����=L3�j�����(�0^rv����8��,����<�Nh��:�@�><2�%|4�t������z��m%Q�75q���k������%�K�(>�i�t��6�����Z�-�I6le($�RԸlT:5`��$�y14LW3����zŊ����Jzs�!�ڭ��i�k`�4 @C�ׄ�F�q-ɼ���T������L���B'���SY�%�m��yT	_'��6v@�~2��=�f��b�j�{�_K�v�D��<�:��y�$?�A��X�6P���;S�V*�mO��u%�9;�
��K$eM �'���\�Q�Rq���8����q�[��N�R��C�^���	�er�6����씌����^љ�
SM�!�p��$�����i��g����7���su5�Lh��`�ϋNsl�`ª��*|c�rfDApˤ:O����G����':;�ٙ��qw�"+B�Er�����l`1>�D&�G?��K��ύ"f��^T��7^̳�Ч�+cm�1�����@�>��?q�u�վvsӊT30����O��c�ׯ---����i �w|��P�bb��7BP˲�佩�.�&����0@F����<,*�\*��x(s`(,�+a��{A�i��0�?#c£��feC��t�%9��� ^�U�p�����N�F����K��]�G	�Ppߘz�Pu.�=ԧ��!L�AX=��6^�b<�o��6UC0Hݣ�]7��X�M]��t��QM���^�n����[�(��n�cY����.���?���׵�BB�%CGG����ոl�JC;�S�N�+�p�ɯ�����[_U�}=���ȃ�(-(�-�"�%����AH7��0�H�Ѓ"9
�C��Đ��{/�|>��{�Aa���9k���>�И#7>j��?��.�V��=���@g��U%,����
�s�o=�l��0ඞ~Y��>'U�褨��L�:&��A&��UC����AP�ZOk�����W���g< 9`�ed�(2�2�a�;|͹�3�2kR��P�S�:X�r��Dl%`�� v��`l�&�����%���J�����rUK�I؅��y8���$n�g��<�V7Z���sO�������b�`ss�>oRhh���Ժ�q\�:���J���n�Ql���K^1�؟�V=F�+�iVr#1���ʅ.|�g:Bŗݰ�\�I+6[S)���,Ze[�@�����L��2�q�2��N��RF�?h�]��!!%����N
C
��t����j���`��� �9|i�+%��:��<�~q���̜x���]uaf�4�}��~��^�R]�~{0�E]7U�[&�cW���
�=#{�� ���S�/Ow��'���M�#��E5r��%z�m�o�7|����{J^y�}j��2";<���g!�5Ri����B�]����5�~�}�w���`�S��j�$@��5d�N\�}���u2�!���r�c.�$�M�,*��=Kj��Y��N������8�C���S�C�$�_|���|[�;�u |�~\�y5"͛&E@.kD��� ���et�qԧ���8�<�*��4��.�9-��O_n�^����꼈�'sz�T�7���(�u@�n���G&C�����GT����4�gw�(|:(�h�E�D�Z��ݨ���'��,U�+b��˵�P7a�}^��Z�Vg3�f�,K�/��>:$��0]_A 봰���3�L���q��?&ߪvb�}�%iDdd��v��v20������%�G���ڧ�{��8�$�VM2�Տ*@�p����$�kFs�cE_pl��z��ʮ�Z/q��M����n�~Lkh�_���7#���6_�L3�3���_�9Û⺖�^g�y\<�1J�ȱ�͚R���ðE��5�3O�#��	�S8�;�ni,f:T���nj���F�տ���mY�n��0�}
�EdPp�H#P?U��X1+	��Nj�o����J��!l1��G�O�^�[w-q떦 �p���C���eB ��k2|����\'�`�b��Oma7?�IS1n?��z��Z;�L	�����W�:��Z!;������N܀���g�`�y'3@&�]�Ε�|�п� [l�X���I!޵ۢ8# �q#���yPD����PR�l��A�]�g ���CCZ��)���V��b�(�ɾQ;�z��Ip�N�J27	����P�� ��ܝ�\���[�C]�>��Đ��~Q�%OѲz#]O"��]#�O��4�Ҭ����8���Xvd��9|�raŜ<@7uT��� ��IQe �"@��^^�xߗ߷���Fl�[d��Ie��k;���}4\��/#��'XR)~ݎ#����� ��K�$���glq�����)s��O�&&&���K��	�G�R����u$}�>�����G�Ć�jg/��b�Y����tjO~4��L��2�S̘������A��c���_9칠W4w���V)N��G*��af��oyj�~���� >��lDo/y��)��dʵR\�=�RNt��S\7��4(Gyf0Q�s��g����n��ٚ�(�i:���v4�qN�0�4��|&6�@L�=ܿ��%r.p䤅@�6v�l\]5�̿�3 ��?�8�չ��;X���^dw�Q�)y�o���=HF�����#|�轸h�[4�fu,��;L��FdB�^��&<�e4(�n�E��T��EJ�3y�����# ���	��w�_3�9�so�DTFXd,�}���ƆNwe�x�%�t�O2�Q���ۮ+?
��M�aDf v;x5ZeE{���=w �xxx ��5g�lp���9�aT� ��M�RQI�Ƈ�r�}����7�u�R��&���C#��)�7A�9�k8� �a㠹޲��m��4I����Su+>a�+3�kʽlɤ����JTt�Nf�0f�-Y��u�bK�a-����UD��
�;��#�Zr�Up�wD��\�D�Y��	S&��,�(U%D����p@2!z���ľ�B�C��x�/]b�֙��j���(#�r;��W�Z��@���1)��<�`�/xGE�߈`O~N�K�Dc�t�h�x�E�J�s��R@���i��n}<�5ģ���"õD�����3�����P�- ��e>�]ls�	�.�+K�5����E~�;�OX����{�%3k4g��!p��Ps�)ǶZk=�����㗤�v$?�"�Q�V�؛rz:y�I���~|��2�W�1�@I����k�"韪P1U<"��>�}߀Td��!��PתN��W�K�F5�1׈*���Pϣ	���EΨ˴�g!�z;J�;�-k��r����dU�v:2U.�ƺ����q	�?D_N�����}A�{ඉɳ�������a��A�A���6����ڟ��7�:^?�lO�T�@�S3Pǚ�|?�^i����.H���z��d�����Tw��;Q�ŖVyt�ȸ�tP��Bz�d��Dl��)b`�iw;�{Q��G�f���UM��nXj]�b�З��dk�I��Y]���X�ks��O����pǖ���7�j�m99� /�ėS��---�� [f�bn;Z%||��Ѝ�x�çCO>U.t`=���<�F�|M��ښi�ҡ�.d���?�҆��r�=�2y�2�+��L:��������Z޺ő"��!�}M��a��\i߱��8n#q�><�����$mjMu��5��]�$�1���z�ćq�~���^Z̿4~7"�����jx/N|�O7ZK��[g�s��=WRx���q�ed�Qo��ۄ[�u���x	ֽ�0PY�ٷ.bT"u+G��`���D&���j�2l|�hT#��s$����l�&��n���T��\����&���K�<������{�������5�nV�17R��A�L�|<��B�y����(Z[\��R��QJB���TRf�6h#>M��mi
v�M2;褋�ܢ��``�A�� 4t�^׻��b�_�6j��q//�-A�M�M��^a�!֪e�3��hh�1���"9J�3��,��7G�R@Gbt,�p�?x�B"�v��Fs��b����G���'����{[�a5OM��1)D���C7KLHh���Sg�T����&�5u'���E���1�����5vI8ť`KK����% \��{#����x��C1�4�����x4z���zc[�J��~dmii�u��ש���*M�[��JѸ��Eqkj�P��Ƀ��x�&nX@2"��p��(._߷�Fjw�� �}�*�3�#�S����5�[��m��ʖ�t/#dc�9u¬7�&��oqKz�X��w�Bۂ��z��� �?�D�ή\ Q��[�9e�U;��η�u�4�T7�aM��9�rU��ر��5g%P�.R�'�|��^���ѡ2��w �^�C�e3*��j�˔�S���V�U����_.�U��sN�zԑ�z�V]�S��sLT4)|Qg<��B�^�l}��y}#ڛ��mGh1��2id���;u2Bϗ.o�Tm�Ib�JJ��ڕ|J�GT�{���z����������_J�#x>08D�����;�~�n�M�$���G�k�I]�S%r��fOn��z��=-��M�s}��娗�]��=Z��#�GmuU%���Q����&]��8��I�@T�;a�i<����K^z#?.�0�S]��/���}��y#���qv���ٝ
V���Vz��då��7@V� 4Fu��)vx/  �՚��������u�%p���V?��u����.���(&��Μ��"������<���ª=Аd�=��[i�j�#/��^��ʅ��;c�@�s���%���d@=��6���S�_��nY/K@/���l�N���s+�*Y*-�l=��H`0��;b_$Ѭ(??hb�Dg&�a��r�mx�PE�7��R�
�7r1>E���LS�q\����.[���5�ky�\��3�����S�X�.�i������V�}j�������'��}S�^��K� �#*d���,���+w��̼E :ⓒ�����k1�����i��'�!��J\�q���k�5�7��:>�\����Fb'v�Vq�p_��y��\c^����閯�K4t���"��V����]F^G>����Ѵ��\�jc�8����������@d�9��V\�~��K�Iۙ;:6���+�v�d��~f�n�P��>*��F�bg��m{��o���q�S�ҳg�9X�ӽ�/\*��g*fϥw<27�G�7���!-���j��M7�^g}*�wP/A�h!
��s-�c�slʕ���1�=`����L_�tp�p�
�_���1k�X����B��&�e��'H�[��y&G T�Ҧ_� �a�ت"A��g2�mX�&o�u�n�����
yq��V�!�x�Y]�'���վ0��a���Q�ҧm�]�	�[��2P��Z"S6t���<��(��@������k����)����͒fyYG�79�� :"���%(e���j��6W�V��A�"[d���?��oj�0�Km�]tlU$ѡ �N���(�bά�;2!l�Ud�l�(���֕ ua�| 5.�� ��s�X��`S*!����������}��H��0=�13��������C���^�0�C��v	�MrLj+��@���w݉���7b&sy�Nt���6I�x�v^DB�A��]��zn���L[�����с5��7��ߊfe8�Zl����g3��O(`�V�)�$(͙7&h�$��j�W��nha`��yO����t����S_�N|N������S��z\���������{���-F�y�b;�� �����P%�4 �[��A>��n1׊�x-�5�N�m��r����Je5ӹ�H�-��.r��Ƀ9�|-UzSe'�����Н�޾=��pP���<"�Xa ���f98|�2�(�`��}¥�ձb��ҍz
(��ru��$�Tu����L��"�Nxnܮ���H���	~o����q���I�u��D�F=�"���-�:�R)h����;zU�w,���l.>C�Wk����wu�@���`�'&V��$�'� �z�4����5;�E�"G7Cͼ	?�9(o8��k�T$�aTE�I���1��7ʫ�6�}4+Zn���9��1��`�;�i^)=�׈���E=~l�Z�@�^�߅4W�:d��G�}+ڬh-��N&� =�v��%s�.��Q��(�#�a�RՁ#>�b�f�s�z�FR���F�	��d��.�)hT�A:�(�bI���W��Ρ��{(**ඬ�/ "���PB���g�U6m�'�&�9pI���r�[�zJmq
�'G��B��̹�F��OrK�W����FB�\�sT�'\�q�-7��4�?��7����c��/�9�=�����h���^+�; �bCC��c{���B�VVW�W��^��V�i�P�5������Q!b��ˠ�ܠ��12x۵'���*ȏw�׭ݤ���Xm��\KO���x���p��B]ʊFG)8[�њ��WA�w｢'�!_�,ڥ�^�V|�v(���ϯ n����-��%�/tV�s�`:E�'��Nm��W^�b��ҥ�����h5����x��|.�j�{ls�V���!S���'Ԥ�ٳ���]����'W����\�.ߗ��4��kZ?C�<�}X���MT�F<k��Yt``��8P �MLL8��S�*j��4���SC�����˕kz#���p���E �0��FT���l�����+�Ic���?�*���a�E;=8J����gAH�҃���݊ļ�(�b��ɷ��n8����P��T��B���<<�b�~(%�%��3�^R��B���3|h������X*��o�׊ �pj%%}��n����0�'��{�k��=ș��D���Bod���Q��Z��L5W|��������P�j�6�CV��'7xF0�cG&�23f�<5�c\w'�@n�3-ND����s���8��F�X��!g��Q�ŵX5M��R|8�S&#k!_II�]����0#���#b�����Ĝ���q��cH�f_I�:2agP��#[��^�9�=2n>W��j�,L�D���稰���:��VC��+Z;�O�%(����ï���{� n}�N���·Cte}�F0Ӂɵ���E�=k@hٙ��������@�`�C����I~�%bZ	�De5�ӳp��j;1�#ur`��)E ���|fR�B�¢����"D7ٛv��G�����f
� ����e�շě�wҬʥ3�h���|�����^ʥ�8�A�Ѧ��K#��.�g��������Z��w�{�����:�l~3Dc���Ԫ�����?ٳRϗ|�0>�^�f�3�^%,�6{Eo%l���5�3������O�b�Xk;;�S=��s��s���zj�Z,��z�v�"r���G�����n�wq
�C<W�B���c��u��H%3i6bHmr-�3�m�j	X�?��4}kB�M��Հ����6�\c���G(�3�A�	����`ُ�0}B��ڌ�ho�^�z@�W�׵җhO��c��g0���>t�3����=�o��ɹ�fn�iTL��ߝ�N���Jn���@ �#p���<�h���Jm'�oǮ4:�X|S���C������iy�Ў�]]mP���!OMF�t��?s����+.=���uB%����:���, 1BY����q�c*=m�M����,G�j�[d���z>-�-��]�\]�3<���񛝀���rmWE_�Z?5Po���%ʷ9�j|6��|��"��ѽ]�z�^P�/����q�x�2kTB}��!��	�H�h�=�b<�Gc'�'2�z�~0�;�0����[���Mm+e�{�u�f�U.=��+;⻟�%2�	8��+++�{~v�2@�u��QO9eU�4e���-�==�6� bv���0�����V�٣2���1`���3i��#H�!���4�Z���6�(����)�֤߽�8���8A2~��~�j�o$<����81FJ:���^"���[kT�����,�����E$hr��A����% 5nL�*$���L�,!G�V��XD:��F썍��6��IW8�Ӣ�H�AB�]�- ��&�Rg��6�0��z�s�M�z����w*.�sk7WD*��t��Qd� }����ȗ��_��H��G�+���׈��@���0��޳�<������j.6]��M_gg��.�����|�ӵ~{��/�ܖ�"*ʌ�V��E!��m���-�7�O��w�&�4܆U�p�0Z��� <�ke�>�i	�,�[��gkF�qRd��]��چw����]�_
lq��90����J�=0^�����^@l�:B���_���a�ɞY�n�Z�"�Z��3��Cm��/����C��
[3��ː���MO��M{{U�O��|3}�t�n �8c�՛�eUo0eB�t��d�NK��A��]�֤�&�1g�x�>��Z@��"�`�hgUT�����Dúz���p`xi@["$(��6i�+)q-��3���;w� Ln���+/�Y��I���{��r��H��5��C<=�Yf&��Z�ͬ�%��{4Wp/��6ƽ�������$Da��a��IBc����5�h������^/O:%R����I`�j���֜��zz�5=9����[2��l��=̔�c���l����d�}�#.�x[`���>P�Ga�l_�#S ����9�
��G�{�*��`E���x�^լgO �	��������nb�Զ��Fм
�f���dԫ�	��Y��"��G�Ɋz���$�Dtj�w�uw�k%�� 3:d���Vy6]�f$�/���o�J$%� )S9��}1((��i�$��߯�t��=�2�XGG^ri;M߬O����[n��a�LTe||�`��zQ���(�S@)� �4��v��Z�u�����'�ydJ���4I��I���1�>{(T���H����q��x��Un_���Mne	�M�k@A��8E�/I�~x�C}>{�,�m��"�X���B<�29(�>@N~~<2y�o��^{e�(||`o_���K�ug?�oT����oHO�	� ��D���iNe�c�`��vuբN�����z��nKG��#M�Բ7"�|�.���t��]g��3؞5�
E��|!#	���ۼS����_s�@r/V&���ܰM����p�u���#+7�՞�(X�`[�㜉�	@�f��!v���q䌺������ވs�=�l�<��5}��Z���'^��6l@�ӏ�ٰk�HX��TT+�x&��Qw����RS���2w�b?�d*�.Հ�Cl��-Y2�{36(��Mzz�?5ï�u$O�[o#� ��� 7Y$z�:6��5P��i��5J
�>���%�
�9I�y�bk �}RNh�G��l4��:��R��e��C/���Pq_p�����i?�����Yu�
T)r9�zl���� נ��������biY�#�UX��R붇���A���D���3򦍒���@���I��X���-+Fߋ2m�/I�U�=��	� ����	���?�r"Nkg�0�Y���l�qR�<�{�%�&oU�f72���Δj�*��* �^8�+����}'e��R<ڮH�ۻ�c��Ѕ��l�ł���o�īh�Ǖ�h���Aq��_�4���r���X�;G�\�v�X+�n�}�$��84
vY��1&X{�t�@�R�!�����~QvK��-����h
�=���C���@K��FPJ�<���BZ׮��_��O��Yԓ�k��c����n֌:4=��hd�O���V<$�äTop{�G���]њ���rp	�������I1���VO���(��bˇ����9�N>�#�k,�w3�6�>&^��p��,�3X��@�;-.m�A��DȚ�$�V��.��PŲkW\��W~�A�庠r�*Q�u��f��Ml�ºE���IV�ʈ�̑Vj���0�3���!��l;S'�ZMS�R���j�OfhV'#���<��}�\�l��m���oC�l�����r�D����+��-%���u�o�~�ݨ���~�Km��ş���=+���>�S�7�b��7��������Nt�[�<�ǵ'�+��/<����P����A�2�X���ȹ����V���?��6��,2�U���r@{"�v��/f����#ã�Y vfZ0�#ER��f��`�qk�<���Kq�� �
^��mju�������׿W�VYw�\�e���Q"�o��E���N��4\�Wt���9e>��&�_�I�N��m��V�wz��7ʓ�w<�g��;q����,�IE84�=ux�I=�����Q���8��|Fl��@�Mg5RH(`�Qe|ʶ����1}�'������C�� sKq���)Ɛ�м9���Hبk�ޭ+���2��;��!�@�m���X�)7�X+��#ރ�T+��-���an}��z:�������ig4���VQC/૩
��+��/��Rq`�O�,k
��6��[�OYk�i�d�e#���ꞻ�͒���&�Z�"p-���!̫�l���&��ZM'� $d$���D�N����w�".8q�Q���
��R2�G�!<#�E�A'"+��ǐ��N�٨��%��L�L��f3A�_��NO��?50�/ӑʢ�lm;��LT��]�̷�5�v�Jس�N��Rc,>*B�=��|ʀ�R�/�-,��j�uZnZ_/�J��`_8l󏊻k�Cu�O��UOJ
��H��j��]�����e>k?
Kih��"Ǵ8���ɅV5�i����o��{��n�>��O*��HР R��BS0�������!���߳ ��)������c���C��-���}�鞵�ؐV
�1H?W�䁶L���i��g����0!���!#ǲ6]dJ���z�n�������٣�$O�Alc{��P���f��vG�����uš����d#�P�
5m�w��h���n�U]���a���k��~�3���Z�N�_���=bE�z����x�WO�8/�� ��l]t�@[ ���T��3Kٯ��.S��<e�������JD�x�������48�uO;��!�?K�{��wn~����PMٓ��*�\��Xx�vR$�kYw��x�J�w�&{w�Dw�(+O�A����>�m��;��q1�j�(��{��B�����(���u�b��Fkc��<�Vhj�P%�z�[/���A���ԋ��!�cLw?׉S,0�6o[8�����n͒<�� �~�.*�?`�q	 +(!�����������>ņ"sg�?e��N-�/��<��}�[^��F�P�3��Tz�T����٠���7"�w�N���ӻvǵ'�i#�GJ�H	���_̳����V;���R��^#��4�0��Y�H�b�vv9GohU�?�7Ɛ;��Ɗ�F��N5��ߨ�sP�/j� �ķa����N4W*��X8t�ޱ�x>�I���m-��	Q�J�={F��i? \��Hrb8p���e���P���`K�� k�[� � o ��[� �g��@aG�^�=OΗ6�&�9V�̼(��/Xb��_�D�:���ݳ��B�hu��{��~>ɷ��2�}e*l�W. h<��/@��4�Q���ރ�耂t�j*�n�L+����n�>y�\�W�j���Pzd�cnsC|�>���:���-���p��'҆`��鷏���_�C;Ya����O,���^ �Wff��Y\��D�PSYlHn��V�C"��A���ډg��:-���:���9�k�ٞ��oj*�k9�	D`K��N=����+�����x��x�:������4$.�iL��_��/&Y�U����S�����F�+������t��6����m)����1��>;�,0�UXRRK"���Y�3y��Φ*��È'�q?ל}�%a���,�}�=]-���YV��D�q�)/� �<
�|:&z ++�Vo��<ǣ�-�p~�����捍O����5�W��i��C͟�X��~��赔T�i�N���s��ϟ��b���䖿'b���'p�@A�.;���:���m,@AS6_�/XY^V�8������ox��o����*+G����Y�C����Fs4��߫�O���{|� ��"�zN8j�#�{�P�����j�}�F����	

�ON��F���,������e��͠<c�a�;+�!��_�� ��௷��L�������\��*+�Am)���{�/�'���If檪�����<�H�spp���w07����5���J4�k��F�YY�v��������������:��NVCqaaH�إ9j���(���Ç��]w0hOmy�����ݯ}����H�,//�.�GB|���e��!|���sT��Q 	�	�����L���3���N����   ����h�hKuh�!~@-�"��\ o	�엿�P�;6V��f@EG�FA(�m��es���('�XCK+$��,p�\�AAA�#kDw���^P��X�&gUK$�SQ\A�����ܯÅ���hmƲ�0��?��r�`[W�8gp��37���C7跞)p�����U�����>���γ\{�H޸[Q��v'��oj����o=��wS��&�������=�n-ߔr���"K�~�bٟO�L����;�s�����W+�@X<�i#��9�P?1�N�cP8�*���6��n�� ��/�q[�l�b�_�]�����<�����54���~����,nթV��X�s[Z�V�+aj��T�<W�S��hv�%���Y.�'P��������L{�m��8ׄ��yDm�/9�\��R6a�E­ixh"��5}k�̰sWcB����f���ס	[�t�Ԥ�%7$�4���4E~���9\�"-L�K�h5u �j��9`�F7&��3|���0��v�ױ��Nv��cw-�����q�I��~Rҕ��I�Q8��v{��_^	��x�BR��{��L�$����8+�����0�u��e%��`�Rp����zn�n�@E��eG)1m�������i\�#��(��6��@q�ݥ��;��R�O�Ȩ�l4E	�ye�]4��1V��Ox��E���m��2y�(	S��FS�� ��-v���,�z�ܠ�H��_$��)� p˅�o�����w����	������b��)"	��E��F).!b�y�]��O�u�=�#>G�);�S��5��:�I��c7d��m���_��η4&{h0���w#B��:l����K��<<<��� }�4srr�z\
�ܘ�:8Jp�LBId-l߭�o��>4��\?��K�$y�����8���P����j��t2~�NG>�Q�"��<�����Ԫ����G>�g ����LjFݳ�f�xC
g:Q���1{@�)Y� ��6��,����Ҭ�x	�h�C?lg�7j
�TNE��8M�9���ic>Z%iT�D}O��J	�9��ތ�]����t%�۷^��K@kxt%�>�
^*���2:
��� �PmD
����|^��b'���se�eR���'�Q������0��Y7��]<He�ڶ��%K�L�T��۟9��ok?	.(ѯ��_x_9���h�a~��-/�V�mޱf`���9���Ƥ�xp��@#-���k���4�Ż�ѿSU��!���R�נQ&լ��\�Y���[���b���{���������+/K˧�ۋ�@� ~�{���3� U.ܭ7�qY��e�M��}���#�����Pb���/��պ��5�4=3<�1�^��E�ZyTKD��Y��k�~E���8Vk�\�dg������
�;GR�"�:���`Q�{��*�v+�w�L�N�����DWJ�4iۭ��j�J�)�1��0�j᧥����~z+��N���KD&rЃs/������R�j1�N�{s��K)>8�Z�g�������q�J'�W!�KB����/��UXN>V<����ɸq��P;�:%I9%�i�˪̓0�����r�G�F���7{5Ggt��n��jH�|{�}O������ ��g7k���4TUo&��^p���U���w�����D������3f�S�)���/�������k�B�;����f�<�=����0�y�3���w*�{�vZ%��������>�\��V?+{��5��򇲘��jhzl-�������2�d{�s����y�uޣ��|���'��q���,Ͱ�f��j-�Ct+�RˢU�����a�Oz�$<���R�ec�9x��0偬c S��e��{_�R�?Yb����I��3�I<=Z�n`Ps*����] #���(��u>��E��zS�{��k�����NSLq�텛�_=��zs����w{��-!!q�8����dk��'��|ƶ�f�e]�b+���)�H���:���է�S=""wF�����[߶��?T��j�4�Y��u%f�o�K�^������<��t��q��[���!S�E�J�\�Ͽ�����/�����n���#�R�ae��fV�BEK+H��ԝ����������0;���['���^%B�ʌ�G���>�j�ϊȬL�ACW����n�wE]��t�nѲq�y���/ɕ�"���wŗkh��EЉ|N	�egUp����@�>�ק�>�����w�Q�8��.wETݵ�]-p(3ߎ�t�?�x����%1�ؽ��;,Ȧ�x��f���u���}+���t�9���o�]�JW����ۙY���tt.(��JQ	a"��Gl�%�a��Y�������+ (�Ɗ��T�]��R�C?�9���|�]�Ue���nz����k�Z�9�S"8`�-�8�%�Y�z�����y�B|f{�M����[�M�{Y�y��9��W�e����h�sAfJ��U�Ϻj���D2�}�޽�A&h_�	
���޽{���VQ'��ic�F���_f�э����O��e;��^��#�Qq�9�)*�V�����C��,�����c3^P�/�
׸跻��dO�Д�u���/ɤ�ۚc�=�6U���5ut����U�H̕D!�ּ5b3ۥf��4i���y��k�ќǜK4�7�`�E����P��mP��fpT%�������	qu#[d^������ <�� ���c���!�xz�������:}���~�ue�y�B�c�h�o��
�g�������r:x���ZvN�7�s�E�()�
���b�����s	������[a�"$O�kT,y���{d1W)�)�Ho�d5ɉ�5���8�ZtZ��mf��[|�w�Ia`�"��;ˮ��'R�m����'�7'������6/�����-�e>���O������P�- 
�jrʿ��^K*:A[cQJʼ��D��2.�JU6�M]QJ5eQ�#-Q�e�Dԉ�e�.o5���;r5�!������W�o.���5\���7���y��$��^dq����ʿ/����*$�ɕ4��ҷ`uu�)��m� ��'���+@���.�+d���DO �	]Ee�*�Yi��G�������i!��r��ȝ]O�Ŝ�����Uei�a�a_��D���d��4d�^a?A�#h�b�$$�]XR"}�i��r��ůA�2S�[oO�������Cg��qF�b��
{��m��:2Sζ�ʻW�V|7���{T���ߺ9S]�#L!�9��-^�*S{�>��j�#����0B���Ĵ�=RW�z�����O������dɾ�������O���,'�f`�g��m�U����{i�����\�x����EB�)���9�Ⱥڋ0�w֯���3�Ĳ\�c�f]f���	�OGy�<���Gh�<R�|��_�ȋ��,���47�ĳ D�@�m�{�}����-�C��ؔeZ��a�'6���ڒ����|Y�x��
Ӭ�| g�"s��j�8�������8O�L��ޕ�������i���iH��8�o��E:��W�#�Yd��&��=ʵ�{�15�I������������ª�5��SM����ݻL�-E�� -�{(y5s��%��zC��y��3����b�Ɠ�V�ד/�k���M�Dڴ�i�ǚ!u�WDu��u	�察
��i�t�����ۻJ��(.��=��
��o�H�(R!7KlR��4�p��t{�ɞ���[ݍ�<�Pվ_��em�f����6"�XD~>��k�9@��prp<24d<"|%�BIy�K��
g�I��~B��`��\���~�eE�U<Պ6����3ۯ�c�'t,V�o˒�|��B�~�v/f@��^�1t�rD�����\ĸIx3Q�����e��?~J�'è.ob�r���kʗ�\��Mk�x�b�@��}�G?L���11ީ�z.��MK��S�`���7��k��K?Wz,-�lnA\;Q�:��O�ͺ������IaJ�;!B��׏~=�m��9�r�p!%(��Af�G�Ї�&�W�'���K>�+ڟ�zPJ&��x��溛�#�Ȳh[E�[]��[�7�i�TxIik���[Vk��$�e�A���Q����̣�o�-]�=蚎f�/�W��~��={4�y0by��(5�ğ{?����}�I(��}�_KfY��0����5�
B^ ��c~>IJ���CH����NM���MY7�yۉx�cj��̄A}�Q�_������!�xJk;�u���%I�R���lH#���D�Y�K]8��f��C�|�9��W��e�v�6����9`L�X��L��h������b �]�	R}��o�6z����U��R���Ϻ���yz�"pv	�H�ߠ�485�ٯ��敤��8xxd��%�^�
��#'�[a/��Ǵj&}y�lS;��L.b��0���sJ�l��FImMO���vI�>0�:G _��-%}�G����'mY)G�9.��;��hM�Ic%��&
T�P��m<5��V�D��d�M�+�
��~"�c����{|�w��,-�Î��[]o)Z����)ۇ�$�<��C{���y�,n�� �R���-��*P��/��ԥl�}���^��տ뤪w�����y�m���W� ��v���j�V�����{!�jg��p�2EE�o%zu�2�
�ߖ��й�"�5���3���ƜI��Y��
j��ݷ�|�N�o�U� ��1�p_;] �������L3��S�Y�)){�m�U�B���1���ju���V�)���?;8���~Z�٠���\@ ��d�����܏��.`�ZV��x���\��_:��k�����jh
�����CoH�Ժ����uh(Y'�pc�顡L/!J�)���5v�����cY"�[�4IS��%�^)��6��3PL��ͼ+ۢ��xP��?��׵���z�1�C0wA��lf":����Đ`��9�QW����S�R��e��9��ش�"�L]P��4�-u��\w�#� L�2��T��$�k}��X���i�Q��9�x�����/�g�-/��wtv>�b�I�#�FcD��B���דfwf��vQa�NS���"������c�=��-�f�
��bX��� 5XP3�	S������w�Λt1U��M6{��NtHH���d�z��8(N]����/p��Z-�.?̇\kT��2,s%#0�i���z���l����N��u�+W(]�ZV羸U'���1S�w��R����xa��]�ОX9b�(L	xz�3-�Z�:���=��u��3v�E�P�^i�|t˥g��>��K_�8>����#����=]|���\��36#������9�����;N�O��X'��,���c��&Ů�	#_�(��;~�A���p�Ж5}���~��1	t<����2!���V��%X%Z�bm�GlIn���b�����ȳ�?N�X�-��k��Sqñ�ۤ����*��:٤�b�Μ%��g�!���B��9o��Q��lR�I����v&����#�0�������΢ϋT��(
����]�'���W�c��� #s3���gq�7�uq�(����wUM�=��'�E��`)���������긨���A�CJ�F%��TJ��;��2�P:F��C���;������?8�}�^뉵�>���\r�z9�g���f���0������,�KU1M�X{^|�k\������~�AL;dTHgb�����/�-1�N+�~�D���R�F��xK�};��ײ�ʰ-3$<��NL�rz~~U4��_3�Kwމ��}~RC���7�w� ��?����k|,�E���	TR��pf��r �K�}EF��wQ-*���F)��lug��K�܍�Yat�
�8�LL��]>�� ���G,�x���߂�Z@�<�4�9��W���]����8�Q��0��I�����U�h�z�؉7`����\=N����M�5Ȳ�]rh��d���PYT]8q qp�:u"���>��N���}3b�|�S����u'giG�&I��Z��}ȵ\��b������C�:���r�����6s�؁'Y�bA�i �6	�Z��W��<���fo.;L89�ޗg�?�yS�b"O�0����'^[WWn�E���j�EB�F�����	~rjhxE �s*rb��2�$k|.��{����b@ԙ�r���ҧ}��`�i��xG�&��#_Q�x������|�B<��Lg՟�Z�����	��8����(����M�)��!�Q��ch�z��:7M�ýp3j<���x��T�����W���+7���j"��f�W��m�W�\7��m7t�����w��Q�k�$�v�7��xY�HA�tW�˨Ev��HCu�[!���#���!��~�+��eE���W�=�j���Q՘+<�9v��9�� $?�N�v)����$���A�����ŷ�&�jq���N�s�^���t�Ղ�z`u�Rp��?�=��S��qU!��{Sj��e�V�k�A�j����#{`��_7�r�هA��ά�l�x&R�7 Х��U���H�pOC����X��t�E��ן_�����F�Z���/���yыɟ�3E�=�����g��������D���rȍ�N�p�}+�3�@�qNif�Ә��k����*��v�"�#�d�!À�+k��@9%��¢����G��� �nǎ��K�%]OҒhܰ]v�ClLI��9�UǪNPd*�!�	f`xo����)��j�ow)�}�0Z������������`�G�DZ_|&���69�`ܖ�c���oԏ����׮� x�ʤ`�����@A��ϱ54�����R��%G#��­�S�FE�A�����'J���b-�a8ڸ����Y@Ff�)ī�{4�.y��|��"iŹR�c��Jm覈�N���ؒ��s W����I9NH�e���=��SW�r`s��?�$�'�Irer.�,��_����IiiQ���ii�i?�p�l�������X���W��!X%o��D��["e2�	e*$��K���w��G��I��e�t��z	BV� -�j[��#*�$��uZ_����0���ݕ�gë5R8�(�UL��j�(�?�I�9�Su?uf_�@6(LT}�����E��op��b�e`���2��q�E�ޱE<@M�5����� �k�|?@��8���<J��ȁI"���D6g`����\&}�W^1���X�&�Wy?��j��I�z��H�����9�T|�y�y<�wVd����Mp�dT��=�!f߬똨
j׈����]������[n�G9�ͣJm�lr@��A)a0�e�Nu��H@���LV����/F)N
�
����բ�8��׾:$��!E,�����Jז�ƺIݯH�����閄�I}�⦷ �t%]���n�dj�%�&���=!�n^9Zʉ���P&��g}�|-K�[�@��+��I�=?l�V�1(g����c`/1�L��󽘰�w�"��WM��1���[DkJ%�$��g
a/P�6�do����b�u�>5�a��*����~T��a�ogs�y�ʖӤ\�@JN�t㐂v�+��ʤ�h���A`�[4�9�M���đY��]�!)����P֠��aϱ�T�4��G��U "���~z�_�`j��@m=����]z��c��;��ǂ�n������)���hh�72��Ѕ< Eы�	�4�{	i��x��$��+����V��*r��K߾�-�'#9�Ÿ�?	������H4����DQ�5���mf5�~�tݶ'n�XiF��N�6�����lR�)I[Z��]���������!*���~W@i�@ �]Pڇ)�'I-�1:Óh��WEK�.i�WZI�>#?�!�"7#x�
l5U?�J�i빬j��2X�{ȟ	���i�N��>���T�a�@
��֓��1��C�T�ꈦ��nZ�y��p�Wt�����C�:�YYh��x���X��$h�d&{�Nqw
�RtZn�|��Mv�UvC�n�"��H�'y��������@S�uJ&�N�[-t_�x"���"S�.U(�݂?-���W)�mn�����������k��s��N������44�`��Gb�L
(M���I�u�'����7�����cn��fD�zVM�"1q�[d��9*�o�dA}T����B������p�nu
�d�*λ�ºո�M��1X�����!��A?���W�kb�&�``Jɝ�M�ZO2Y��'����[j��]���>]�m?Lz.��&N�*j����Un?+�]�Y�BD��?���O��X�u����2�ֵ3ړ����}��ʔ<�����`P��q�q?M���)"�G>���9�}��$L����(��Rz������7?Yp��cp��C��`�J�`'*K��&|���|9�Wd���ٽ��{���]�C܊�Q(�e�ζ'�M~0������:ܐ7��IL^^�\S�����8�Z�Q��F}����i)�p��qkLfe{�g!��sf�tA�D#�g�z<��#���b�u�6�4��%%����� '�c�ꍠa�}�@{��^�D1G,��H0��a(	�Ltr!�s�z��*��"$�c8��I�'&<�H���iC�iC�������f��g��j��\l-��YiC_l�=P�FSt�P��f���	��f�!�\o�����ˑ�p���B�w����bl&��VT���\6�\�����_3O6(ZM���K~��+-�P�C��g�|itK���^��z���Mw0ڼ4��O]�O����Ǔ��� |�Њ��E�I+���9�����eZ�W�­���V��琏�T3tќP2�Z�;o?�����5�D|��̀��#��Z�\�pp�0�"`�H@����RP�������W�����e �jz�$��!Dt��X��e������������>��:n. =Yax��� �����n~�P7=,����p̄oU����� �?�#v�?����x�S�K��ǌ�O���{�P���W��|哺&VO��:{"�s5i_��^8����s}�H)i�p��1��Ƅ���n�1��^��������ff�O��%�� Ҙ_��)���V���Mzv.�Yh��,���}j	
�Nͼ$��)��^�qM�Ɯq��<��-���*>HbV
�^A���잻�D�b)�I�8�! i�X������s�,��h��}ʸ:��`�b��W�n��>`�λ�x�8F}0ܫ��Gy[Y��Fs9y�-6�d��@��t7I"lDB�0k�
���E�Y��;[�&�3�m���/�0������=LǱ󢹚S
O��C�'UE<َe>��F���UVr� !��t��wT�l�-�X�1��sd��Ao�MG�X!��r;��le�&�3]����-��&:9c�jD���Yfi�U��B�r�%����o��K���^Hym/࿖��� 5yZ����L<�Mt�h:f�xh�U����>�ӣ��]���Gz2����8���;T:�j>����Z��ޫ���

n8�gffTc�g�M r�9`j�/5�*�;g��,�^������%�n��#ב���Yg�4�f�]���\@��}������w����F��9d��ĉ
q�����B��ɤ6/2O�@:�U?���I�4in}��0P^�S�����/��/��G��Y��+��~��ZΥN�A�X�Q�˦��]*@�s�o-��וNYqd�sAE~Rh6��i͚�HO6z=K��p�d����v�(�US���2qܷ����Mw�a��O��g��j �/p�4H�7��d�Q���r�l��Zo�_�'��v3� ��m�@�4x�"b����j��<6qr"r��~�U��PGZ8[�N��4a��P �� �Y�#�� �n�֮��Zg�����|>�~��q�7z2�d(��EĆ�+c�{�ړ5=�'�Q�9�3I�w����-Tb�=!�x��ĸ����s��w��-hmܤԇO�~a�Ff�&6-�D�(��"�t�m�wc/�2jj���^6���y�G�dq�po�+
 j~�q��T6F�=�(āÞ�!�g8�O6����I��c��_�0�L�Lz�X�˲J�[�e���2\M���aք����Өyt6�6�Ǥ�[i��c8�j�(0��x�@~6�M�2�}Q����hJ�ƺA�xĊU����@l�θ1���g_sG�UMaPq��s��v�S��G� +�]�/o�6w-��/�l�|߲?CJ�4�}w*����n�C=Oy����eZ]_0呐�;c�Vz!d	B��Xfn���3RyY� ؗ��a�/��{֜�fu�%�F,���Ђl�I���;3��	��~��������М$0���W�Y@�sB���rcst)}X���W0�����s,ʯ�䤄��# 8�
�����췳�J^�7�2X���!V��Y�mͶ�v���X;: Y�����a�떵P>����<{{��e:"ޯ�'~�
�	I��K����zڳ+T[<]y��r�G�5���D^:F�t�40	�0k���'WK.���)��;L_�J��=K`Qz �J��ڃ��
����xA5��r�Skv1�����bԇ?�v��IW̄�*eq�����tw�b}Y��S�o �_���]?��}g���@H����{��A`B�	�}�S���L�K���
�"�����{�����R=Yr����ԡWoP)�Q����/�Z��.�ݲx���HB�%
�@��؍%E��ӄͷ�.Jc �����X�|�vy���w�r�a��c8����y�&~/��l�7u'�S]*�%_���MrK���p�r�zLe&z�Dׯ'���Y��=.))���j錦6��A�� $	8��;�!`����=��v�`}j��J�|��q_Dla�r����s��P�Px�ڸ��#�s�e�:�{%#�	y
�mnd��GYD�Dhm_{ٞ�9���<0k�J��M�)j�M��`�\�����e��HA}�'
��ĺ�2xhN4W=���C�H��@�����Ty?,o=-�h�����+�vY�����-�8���ҊT
���Y��G�����Dj�/����?��őI\�g����?���&���ؗ���X�/�vP��u2����*�;&�xx#�� ��c�S,i�R���-�o^�n[CY% U�S����WYm�=o5��
���-�Ơ�B���3<ե��ԝr�Hf���������*n��M�1nv�*c�K_ˌ`�~jީ�#Eޡ�4�ƽy�����t�C̥�c���5�L��z�C�;l�7v)�n��&�վ�_�w� ��(O�0P��P�h@�0B�o#��*9-8��1�F��
��l�ʘ�5m��un��Fϯ� �,��K� ~l�C��[�?[VxL��n��q/,����x���~���!��4����aW�:�Ô�v�����X�� `a���-*��Uo�? 4H��Tr~m�h��v&>ea�b�-��3�fF�F����Z�XV�2O�F�Q����,<> L��	�o@�&�'/��6��S��a��Ao�>��6O���oH��І�W��o:β�x:>��Q�>�
d�4�d�!$6'����䏌�G+��K�h�?\}Ǘ�i���PU�H.۵�����>;/z,�|�	�V#
��=��M��a(B�q?u��((��Z>ʫ����/�3?%��,+{�T��9�1�q�.@��{aa�����@�2�"��uCY_Ai@j�������=��z�!<��4l#/T$��}�^�k�ͣ:W.ÇJjo?G��b�=Z�>���/=nWv>(�p�e��R"�#��O��\i�E��*d���5M�q~��0�����o��̪}O����MTQ�w�t�L2ϛ���Ƴ�]DٲR��H*u�U���D�Kl��P'���+���鎔L�N2 ��Q�_���I��%~�=��L3���--4��9���GAA0�?O ����t5�k;��G�qTK��^�k����b>Sܥ� ���2s�e_��Gw[qrr��oO9��I|6���P#��B��!���{cc��h��"��o�^L�!�1�x�6��P�r-�nʭ��/�^Rs��`0��.=8@빴((�~\��IVE�\�ͳ�/���eƸ�^<�n*3��ڏ/
޹64H���d#�"Sw���w��p}`=�^v4c��/lohWRP2E��W`�T^�c��D�?�`�.���]�=�g��48f�����S༂td*�|;�!�s�ykp���M���=�[��"F)�l����"��8�@��*�i�u67��5�t�.�}���8$DK���#kv1�	b����GKB��~�mg���&��A��csF~*	@,cOj���L �?��Tʡa�+Vz(h���o����r���Aj�����>��M����R�_��^E͑[Jy!N	*;Jd���	�`+� ������3�_�w��ޑ��eH���hc�� 	���Gi9�&b���WN/�j}��Z�����SJJd��u��#��ih�/
�5���o�\s�)��]��7O�Qx�l�>��{�>y��hn�@��؂��?����w!N�~+��F	0��d��<Q~x��n/�  �Il��
'�6,t#���O��HQiF��yA���p����T��SC�����P1�M3��cG���V2�q����/�w�FffzQ�:��ӭ1�x���[IJL���H��A�ݠ�̴�Pt��x)�x�9���E;�_�����#ޑ�^�; �$�!� ]�f�1����{nM�♊�#pQ�P�Z�3�o�Ҕɘu'�a��[�X�B�qǟ���v�~��B�T#��E=E�i�:��� �/`�|_�#���6�>�����(1_c�F 6���2c��vؼ`nnO�p��&��r��\X!`�޾���C�hϠ� �\���l�^�GIt�|.66p�;�x+鳕�:V��ĕj�	�b���9o����ﰠ��޸
0/�k���U�0Y%粦m��dT��Q���N>��;�J�ME�+�}���ո�S�/ՂJI�h{�������t�����J�x��G؆On�����ҟ��\Y�}���/��NvZY���cTv!GrJ���|tY�5.E$F|��)q��{���o�p$�C��	��Ce��̻W�;t)���D��1��ґ:>߄W̖����٭��I^��U���!�_����D�d��.�]U��Za�5� ���H�l4Тk� ��/���4N�tA����U^G�h���D�_�T��,��(��;�3��O�1�"Re��H�nn�����a��:�TY������=�_��z0��YT~C��<�8~OFN�w?�s�� ��}.�b_��]�hǃ����5��ZD<��!�l���WUx+�t�Hp��D�̌[�#<��L�5�����>X��WJ.d<�[� ?���TÆ4Ṃ3f��^؅}�B��F�t�[o�ܾ��:aQ�)>Ⱦ̜�Nyſ/4�A��q4g��,f�P�ł�# IL˿�.�<33��w�hKۅ�/�(HJ�l���$��͇�8o/:���S4�`'*}�sWlY�!!�����o*�z΄IO
��-L�U���kBQ���Rۦ�� %U\��U�������J����q�_�����A��0��"���tdc_�=	5l�	<��Pa�h���Ât�b8��>�/�2z���9XM����e����Q���v��M���L.d�@=����4`�⮮}iG/E�5����-S�/�� ��h��W�v���H�\ �)a_�9�7<W4
83���;:�]���P޿A� f��ޙ���`N�瀩�lo� �����[�lPb��$���-�����!qbbZ$�ߔ �{�v�,I��#& ��#e��d .��]m���FȄ����z������/1�G
@d4��3 �(�D5}wq�SE����PJ`DG}� ܼAl�`G��/����!Nv��pynv~��ذ�}���gn�Sl2?-oO�YAgO��PP��c�z1��Y���N��A�~˯C_���&�?=1rh?��"�H����]���v�FOM�L�\���_�~5o��E��=����̢�!��My4 P��ֱ�$��3݈�B��"��O6�<jڧ;0ѣLv���9�qC����+ki��I,U�~�ϡ�6U�ܗ5����Exݵ���V��]?U0J@5��d��;J=��:���k/��M�<`?*Cd�,�k�$0z>�b�D��]*k⽃�" d8)�!���!�C5X��<'V�����n�,��f�BQ���0�~�����H���=uAzJвnXzŴ|�c��p*�)>�_��.׾�Che�r�v���Tl�kx�<� ��f�s/�Ũ�3C�ݾ��ւE�+gt8{A�R�h�*It(i���$�1}��xm@ʇ����V,����>�.@eL"O\���F�s�8!>��ϜzDѲG�Ee �T�S�������^���wo�d���=?DF�})i=����J�y��N{�������u�_������V؝#�iC*���B���Kvq������.lǨ/x�_7@Vg�j��tP��s��p�/_����M��О�܍G�K���1��ė
��5�� �J�'Z���?ܽ�4�׽G�lx���A%)ˏ��U��H�9���W�G�.rh���9��>�9�� 8�ǡ���b�Ε�D���c[
Hvܛ�.��%�U�����{<^:o0�����y1�����W��	�>����ͼ���6�-l��5����;6��6�U�D@7r�X4�ڪi��M�
CV ����?s�ܖZ�qFܻ���d���`#�(��Ξ^Y �~�#�@�q�#��X*R�AǞ1�D�^Ķα�eP���@�cf&�Q�D���.V��`�;�E������'~�b��ܗm�����'�o�^��I��yx�*���Ȕ���=�ѳ�}����Q'����j۳gP&��\�,?TC���V�RL���+@�d���-�\�_u��T���*S�w�6�it���Y�~d�^�?g�5����}��o�ɼ�p^�rm������;P�f| ��0���i�D���qr�m|���?�1�;	ĻRMÙ��3���XU�s���J�������Q�ß���ˡΨ�1��H�����1�5��a�jN��F)���7�,5GJD�k�d����
  �a�t��V��.��CS�zrb��X�~d[�3
 .��<T�(

#J�jL���ۨ�ԕ�04��G��w� سl�qzIS�w�٠�r�S���	��M�
}������R�{3�hf��[:���������h�^��������0B��̒7]�}Z�bM-�K���l�9�#��G�O�%�Mm��]�_$n��1��.���:f����:kj>���{U��\�vmg�I�U�ؑZ���ğ�<�6 ��k���DOk�#(�;F�] 	�:����Z�9kK(��c3-��|@��5=��i�Wm]� p�V:�?�?�����f�G~>6�E��]e6����B\�)���b��\�Q��k���t��X�k��'�	��� n��&�&~2u(O�+9���&�qQ�����g�kJ~|�s
��2�VLf�ש�֒�ƥ�����Y�?S��B��G���F-#��X;��~7O�T�7�d)�����[���o��C���
!ɱXv�љ�!I�J�a�񵄀�L�Э�;&�	�"Jw�g\���b������I�ܴ���vX��Kg�&U�̇,�{Q�lN�Ԍ�X��{�=�kx8O4�d�/$%Z}���4�a+���]���|@:D��<� e������z���:�2�=!��S�co��|&SO�+�
����XUmrhSu�����.A�6FDhA�A���"e1�OgwZ_"
�3p�\d��|�_�/�8*��_���J݋�2K�%{a���8��v�u�[��`&�/E����\���;u`�e�r(�\�-�(����op�l�{x˪���O��q�,�����x�*[���_��������C�:��()P�^����~�h �>	
��C*�)k,��Z8�l+C����ijIk���k�=@��K�ay�C =P�=nX��2vc����,��@X&u^j�r����"���G�x=���>F�,s�&�����RAC��U�Y����B�%�{��P�D�q#X��g��SN=����u��8q������������y�\Ũ�W�e��U��'��o	@�ii�:���xD:k��[	�<�#��}h�Wx+�-�=?�v�L����(���3�� �hI`��D���?s�F�u������k���{ܔRa���$,�t�}�K�k���ʱ�$A@�V��D��� ����q�.�|jJs-}�����M�K狡���2uO�ߓl�FT) �Qr�6�\��v��� f�C���!���˩%�0��`rKd�I�;���e�����)�,�u#k�q6���w.ϸ(�dp�wR<�v�s� X"���#��Г��� �4�HR?$�[HH
ֲ�*��o.,*I�eV6KO��t��.���ELdU{@�2�i�.$�ԝ��B���t�����=��˨}Vz&u�1�J�Kª~��w8<�E� ���w����E5
1-��E,�bt�OY���۴�lAV`L1�G��X�֏{c��P}�5�hՊXOZ_s��Kql��
�5`s4�9��&���_�j����)��ȃ:�Y�꽪��R� G��G���L��'���Ş]��=N�:�}~�%g��%9=҅�96.s.�E��8��i�E�[�Z����?���7�5���g	c كȡ� ��䀿;�%�S��gR��y;��!��WOY��:�7����\o+NY�����LU���ݫ�_�&���[���c���������N6��TY`�3����
HL8���P��{t,�-��w�-�/����~~N�YO�T�j},eϹ�s��,̋�]�}��7���;���]���P�m�s'H�{#�����1�?bEz�xCrp�ܰ�d=~D�qc�UW��=*�*�s5��/T����m\�x?C��/�a�f���d;��N �x����.	u�n &�DIm�wCɪ�F߸("M�r����~��!�����:��
G-D1�I�r�4�xJ�OH�2�Q�b��ț��[��=q�
$@��^�' av�o��L�+Lw��=��;ob�	#e*"7�����P���]-�*����?�(��2�ÛH��B��X-]}��&dt��$� ���a9$�w����Q���-��`�����H4��~��X;�fߕ���Ͷ�"^kR���m��o'U�%��W�Y�RЛ9�}�:�3ts���mbI��J��N��,���⇉]*>�q_��x�G�3�����̻=�<�f�gÉ�G3����_ �'�E|�ך̜oL�� Xĭ�zE3[.���E0��F��S�ʉ_�	PCX�*�D�\������y�6����)�c�2xKK�ZW�����?��D�����g�g"��G�o�,6��d����.(���:�Dv���z����Q�1n�N��|�¥�p ƌ��]�ݫ��h-�z���wɳm��>[W�w����,��#~=��p�L�sO���9��&Ou-�v�"�_m����MO�+Bz:-�P� 3}Y�t���Fy֝3Ӂd��
s<&���䐲��p�%���=�W��m�1c��LQ�R3�I ��F�\��G�@þS_#Q��Tx ��_DY��`�ϣ�ܯ3�\K����rp��w��ڡ�A��f�B��"��C��NI�����'U�ETӘ�Bȱe-?��Xe\�h����_	�Ӂ��\B�7���a'���T�JFT_�^\��T�/�LK�yJ��k+d����׿�b��w�/�y��Hۦ�-�zh;��%���˽I�0a�β�Zbn����h���O0v��PO�Ǵ�(d���,� �#�,�=&�օgZnUZ7�&#O%0��vHd%|��y�"mC|h<���������l��L��y�-���\���aIr~���$ �6��<���}�f��=���g�Ge&�?&:��:�2Gd�$ �O����.�]��3��U���#ZǢ��K��/N��u�������Yȭز�7���Xb{B��^ƣL9��Y����S��$Pi���ا��� P������{-*����Y�>��6���A�P�x��b�5�u��Z�%A-Kۉ�hSb���&7d�s�.Cz��&E�3s��c{FU�Љ��ӜR����ʅ�嘮^��)��=�C�7���M�p��!��@�B�3�e�S$��������j�z~�뒋&���w�Og��rLty���@�/������0�|��]�d�F_"�@ Քή.~~�##j�w�c��U����W;.����g��t�#I�����H����]a���m���5ɷ�j]�%���r���Xي�aݱ릚*K�y��4=�gT�QZ�z����CQ}@���FA��5��7L
x�M��,Ӌ�}��
��y9�oM�͊[W1�M��Xt J��z�Mb�D�Нb��w�|��+�����[ZM</&��9��K[�ﬕi�k�3�@�<ϟ�������t{�v�� 8ޙ&�&��'.X�E���X�..�,\�������C�RF
���.���JT�����_K��Efa�vn��]�Y&	�<�TP��*��o�2�䚲[ۧ
�4ez2����׎���c��-9ju��.Ksr�n��	��O�X~ֿ�]���5���Q\�_Z<)��C��M�5׎>�������T���\PpMҽ>�, �����n����= �{&�3ms��i���ީ�����P�1>�Y����=�Y3Wa:;7��j�
& � 9��۽��@��0�7e��|�-ߥ4!��z܄�˥G��%&��k]���6Ƈf��9�-ebK㖶D~i�.&��</��.�b�1Eag��^�<����&i=W]���)�z��SC��F*L��9V�CQ��5e��3��^^l�����CB��b2���A��q��Y���hť�3Z3���$Ҋ��EӔm��TKw��G�U[_���h�?< E����OMT�=a�{�ލ4e���Φ�����*��79~'�ɾ�u�uw�"gZ~��g�kVS��y~����J�	�i½�9g�l%�-�]6_��#���24��-&*M�*�~��vrۮ{!�kv�(�V'�t
j�&f	���T�����Jƺ(��20��1_";e#��<��ӶL�̎�$����pՑ�R5���	�˂D���,v�4��Y+eoD�%�?]}�����{�z�<�%n�@��6��_YY��O��6��9�]��He�������f����������~[��_�J�	F�e��ʂ�����u@�{�3�J�T�M<��c����
������.���ELQŎ�W'��F��E�➃���E�ye����ޓ#����ː4k���?��!�>�Cv��.xk�����(k�O�=�7'E��
��8:��mV���0���,��ty.�TX�������ڰ��.Ὧ�z�V3������1�axU%	&�ጴ;:�I��+�q���dv���,���x⃪z��;�xFT���8 JT������ǞQs*�/��q���bh��;��r��k7-hЄ*�}w*
Q�Y�i���\�<�.���{�nk	�G�D�a��y��7��g!Ce��'�׍�2������J`�;,�}�P��.Z�=�����gz�#$P��o�;��^�;z?Ú"�ȉ�����8��j����㘥��,ˋ��{�O��𬋛�n�|����I�w��1K1�����,�{��4�ǧ/)Ws��7��[%����H6��{~�H����6��y�~�$�-%�l+녧�*�j�y�����uܻA6&��<Έn ��Nr~Ì��f��};����-�P��s2�04�0N�V���#e�6��G�ͺ��T�R��@��%5������4� �����$����!ͫ�����	���^7�-֖�������x� Dns�,�Q���[�HF��
_>/X���wR[�,e����t�S�ە)[!���j���<����,v*�8x�?�S^����m��]dRz<�0��-M�xV���}9,7q�~���� �X�!"��y�i��!�[^��'R�KT�N�	��r��%Z��TIyM��7~����e�ۛ���>n��+��5�p������2	a�����-�wN7��x�c��N�J.�|r�>)`M�ů���~i#U�Ej�Xׁ�󹂦�^����<i���E�o8`�2��S��d��O10�r�5��)��2æZo+��DŞ4T�w=��2J��Z��qh"���lJ�6����`�U2��q�Z�nT�ө����-���(O����~�ѧ�u���U�JaM�V�F��]=F��F��8��(7���3��g�K���̴;ߦ�.����L{d�'�R՜k��߹�ۿ���:��ƺ��_/ݤP�~t`�B��ǉ��tغ�9q�[h>yg�����z��L�`�ۿ���xo�~��)��tn�A����~�)a��ӕ��	wC��ߕQ�ǆj3�g��g������rԻ��/�4R���]rG[�{'��`�o�V��w魮��P��}����e���ϳ�*�\�oORW[G/��c?B4_e���]��;����rO+�Y*����DU��O���i���v8��<�\{�w�oFԚ�]����KƪQ(��p�6�@��fi��բ�gR{;�˥ Ih�������wu�������&A�bw[*E?~Ȕ��:�,�����l�ٛ��)7�oc�ﳨ����v*�8a��)�9aI%���?>�(qv?�|[Ԃfάk�aJ�[����~�cN�.�p��j��۫g�N?d.�a��B�*kYL�n6�9�(j5���_(�*MJ�� @w�i����,��Z�C��G��	��H�N�#Dab�g?J�,⯱�������n��ߎ��kԬ�Vq�����y~��U]<�8��qh�m�CQ M�3/(FG/�"�E�����C���޾j��`^���n��.��Eo#�	Zs�����~݁!q%.sG�+�; ��|S��������)��������L/SȒ�zF5{\��{(�i$5sT����ϰ ���F�K�_�t�����y󅦁�b	ϛY�{?��:{Rk�Pl�
x$�P���Pԣ^q۪2($K��d�]���H�"KBrr�Y�(������g�M�h|����&��N?m�����r��Q$���,<t ��dri��j�2H=P�\.���p�F�C��QLa3�*�q�����d��h +�3��^�y�r1l_��V{<�{X�����_�e����b7D�i���J��-�ꎌ_Zyف_�����Ny�"�u�8#J���T�����P���A��m�[��At�i6� 5����hV�>+_��d��TV�ta�3��l�
w�i<;���7В���v�@�lP�ca![������Pԭ�UY���G�9�zF�~�6��w����MCS&�̢ÖC�v��-�
�q��_���a�c���;$u2YP- OA��q^)Y�a���~��/�$F�^*�fNW�Թ��yL��`������gy[�7���b�|DJVwĥ��)����j�Q<MuJ5�l�R#�:%�6���˩ʦy��N��� ���~PL��� ���{qr%V�ty�D��N0י���233�i��7�R4����L���vb�I�Ǌ� �Xی4�=Lq��SZi}$c�'Z�9jc�I%̃g&���΁��tM1�v���RwB~-�xWw���]9��$�l��W���1>|m�r�6$z���c�q��!��m������Lԝ���	�s0�Aj;�
���o7�ĕ ԒGj*8ǵ�Y�xN|ʧ�4�P$ A�?�&Q�S��i�GT�5Zנ���r�h`�3�`�Xڱ�;hm�.��B���������j�U�_���?����SG,��vvz�Y�E7�%~�\�W���*�a��x�%
��=�e�E��˦҇6�Ň�ch����w��+�o�k@d��T�(1�!�F��ơ�����eM�}/�x���)ۧ�}ȣ�4�`�3M�U�Qȷ�̼���/0���e���|��bs�G
�Ozc��cʏ)T$䋕u͜qs�}����8[��nb��ܴ	���⾨���ۻ�l�R�=N���gq�R�o��/���'YrRD&�� �@���>y�4��(u�l�Ѕ�t`%�y��P��@�@
��x5�-\�?�:������>��հ׺G~��z;�_��QM}�]c��C�����������H�tK#%�%�)Jw#� - �HIIw��t	�P�C��9���/��}w��r��gf���~��9��xA��q*~�c�;�nVa#����j�M7^ͺf�3�>�|�)-
��}��#�[���9�)����<c�J����R1Y�rT]fr8ȈI��W��(�=��hHIK[j#��HO̤��������á�����ѹ.��_w�3�ԉ�;E��d�5��qw(�h��4z������_�	;�� 1xG��k=�H��']�G{�ښ_��a�;����֥g@��t!�'�s~Z�&�,/%�;ߘ  �y&�gN����V���3.�
����h�B�V�����{8��a ���&���7��
W��e��k��;}����nJ$����d�x]�z�T���߂�|�����t�Uhc]��#����!BLC���5�b�s��:,n7�b�
8��J��K$��U��G��Y���m��o�ϻ�srp��9��C��=,�1nC��W����aþe߹3g����~�h�������ɛl��O�}�[	x�W%y�4�J�D;hƆ�0�Ϗ ��/�v$����$�����9��贁g�4����v���`�������f1��"��#/�L}�Sax��έ�+KK�m�sk��є�"�N#N��5;�v�
s��szgL�^�(�l�В�}�dlde"P�hl��R����'Y���;m����'{׉S�|��@�3�f�]+V"��l��!�`�ި��-��6��؍�։U;�By�Uc �3Ky���<�w��������W6�M��C+g��w�M��o�����#đ8x�P9"��P�W��L�É��+���Z�����o�#����b$�!S�L�Y㤁:��=�y�dO�N�+�jmqmw�r�� ���r���V=3`)�ؤ�3S�e\�X���,k<=�+��
\HMD���^nx��ާ����gO�p��D��h,�?x	�-�O�(ӭ��Fl�<�Ck�e>�Eg_	��e�S,�E>g��D�
*��[����pEy%�JG~�
*�2L%��;ڟ� V�CgFd���l�Z�>�c�&��-�T����8�T�$;�(иs��Q���7KK�[��h�M�{�
�hl��!z/��.���2��Vtfn��IC( 3�,͛������O^��n$�c6�� *6���������U��k��r�#rک>J�]�>�����b%�yK++0O�x�C�;��S;�6 v��|�J�?H̿o�x>���mi��q<{�;1+<K�"Z������^:-�q;|1+���j�����+����\C�dGQ��Uζ��ӵ�<�ZN>�$��og��"�~ڋ&��Jc�y�g�g���
�L����ʰc�{�7'��-Խ:S�:F�C�%���V�o8.n�5$v7�uZL�3������k�����8�|��733������tW���P�%)(��o���Zʒ�λ��ٌt[m���n�=�ZW��10�&R�Y}�a�jA��Ӹ�0�1y~�N�
�۰o~ ֧1��=����@�!"c���mc����G�.����Kg)���鬮���&A�Xs�R��f�O�s@[�4����wh�_�ȴ�uձf
P�H��(J���z�f�k$(����<8<��Y98� �6�\����c���	C��C���!���i��_�"~�%py��s@�[��G��
�}����8����'�u�O�(
]&��`��h[��+�;��uO ��DD���H.��w�"5=�
P���؜���e:��K�\U0C�.'�F21&ڠ�Jw3lf�ݦ��:e�N�������D8S��;���D�(m��@����xؚ(��\���#s@�͍�DK7���N#^�B���H XA*�ٗ0����%�������� '3�	4������� DX���#��7�W� Z��Y[N�I}/��u<�E	3�Wk���|�Qic�Lx�B,Kt�2N�]����`K�쿹)80D6 Wz��Z����;�����h�Fɴ�Ƿꞔ��LU�E���Ȕ1`���2@�[�����s����vfV�����u�`b>deQx/1�0��P�Qh'�-��,\6��/�텓�LC�j��Y� ��	�yW=�hϗE+��1RRR����s��e�z����%RG m���Y�6"�h��%�w����jq`` ��=����.�]�����1dLҸPaξi�d�<R|#?��C� J}�'%��[S�̺5z����yMؓQ��2��kdf*����M,�[n�w��!h5Ba��,Y�n~���EӬϹ�Ҿ;]g�9g�>`D&d�|l�B����Gd�W"�;V���OSӸޥ[Ih"9�]c���@QFk����W���t����9{N"�=i�q~���/-a���t)���[��� ������V���w�������I䂹��*��'!*������;(��U�Yz[8�'�#j5�K���Oc�ܹs���-C�[������f�}%�a���D{�=qő��L����A��L6�Q�Qb:rcI�#;��Ye�sq�==��7;��ҷc����_�d�:�id�,�1z9�e�9���!������r�K��N�ʐֆ}Q���s��m�OG���!��;l/oo�������� b�rP��=ز��U:5�P_V���� ���Z��$�y��"@*��P�͝�ƀ�f#�v�׀��������˧��GT�+�r��zL׮9W��Jf�ѭ�[��y�	=9�z�EJ�J�g���jz}�E˘؋���O
D��<�*�o*����-����Kl1�w��nNHA^�i����獭#���{�d3�tI�om�
�nYmMU?h ����W찈�:�%H�E��7CԐ�]�@�X���@GC[�Q��Қ���������R����p�>���֑��h�e-��,^t:R���
�%~H�����I1O������zQ������_��{��ť��פ��[�bF�K��:k�|!{0N�yW�� ��_3Ύj��2�U�W�ˍ�ww2P=ަ ƒՍ��Yk����H�هd�k��}]p�QeIDu�R���������$!!IIJ��������ZH��>o$�n�4�ΨaMFH8��$��!��k�㓮�ׁ��9[7���Ҋ"@`��&Pz�r"�=ߨͥGRן4�����M�V_
kk5��X��<}-B�\����K0�`��tO��c��T��a^x�W���]�r0eUF��O6fye���� L:!���Jˇ
0�yW��7�C��UKݗ]�\#����z�6�]aR9��f��C-��q=��2g�Z^vEƗ��<�����~6744��n8ZT��0w�䞞��1;���v�P��ǳx����Aن��������ihm�[��C4�!pf���r��Ƹ���;%����@;[?)�������l�D�gz��e�Z$�� ����d�Jr^!@L��ƛk��˔<�,�5�	���+岦�a^�kѣ� [�1��P�Js��1��"2 �WqR��`��̟�e`��ow$�΂c i22nf�I�~=P���4�2�z�~*(wdo�������&��J��D(�\?|��A��S��jA���{

����A��.�ߓ3��lc��8��������=$TB<6�!����A먶����x���4DGGǘ�NQ="�G5�#�9ZL���@���°�#TTTB��^o\�u���R ��Ϝ5/0Ho��lN�}���v
�4�1춎>��@l�%�7���/��R4/%�ۥFVx-��qN����ùh`_@AA �cI�B�	DP5��U��+C�xg�R�$ײS�¯l
h%�*� �ڐ4�� ��6&���ނK��Gn�����<o	f����qU���=pam\/��e\�/[x-�VĜ_/���� �MO��<�].�q�p6
�Ӈ��9p>vZ��N0" 20�G� ��~�Qw��p;WL�b>H>���_�6=ƪ]�$Ϟ�#��Vh�Aܪ#�%�8<~Kt�,�t7���夤��&0��Jp��}&�x
��P�ܥ�v��f���*��0�F����yˬ׾���ӷ��j A�ٳG��=�!�\ 	�r�:�icIc+��9�~q�t�kp!�3!H O�O��7�}%���?�����6{\�ϕ�mbd�x����2�N��4�`���^�ƣ�y��<�A��A�G���2]ƙq�q*��OX�i`���Q���/e57$����
�7��GGG�j�'���MsU齏��6�ZK1}O:tZ}�?d�
l�D
��r�|��G2$/4O�
��O��#/�2���MMiT2�������0�@42�b�8���r���֮�0���|lb�Qo��ف���nG�V��5��H__;�x��Ӗ��D��O3ė����>�&��T�\�|����t�taB��7N�ԓ���nٱ26�XXX��}<<<�[�v��^�Fؚ����7�m��~9l(����"5�)hg��.�G�Z[�0ܾq���c�p��ȍ�;o�i
�yy�\j��"�~���ҽ���f5����Lz�e��Wz�O[�vD���d�8��~�ꒃ��q

꯱A�d��8��3` #��TٓGݏ���*�B?�d���2w�ϥ��nb����bn���[Pyp����~`��@�ǟ�Q�8�яQd���n''���������<��;����#�BDܲ���uZ?�88rV2|�#�����yy�� bC6��Ah�Q7˄�bE�����9�Lש����|�n���M5U�C�+zxx(�󰡱��r��(��[E����S�?�p��fJ���Gvw?�9�JK��:�z@��I�����;^��٫!���Jd�&-Lman�T\\jn�����êh�)y^s� ��^[���YÅX����zY[���+�yGtӫWZ��œ�R�	\������8~x�
���e�Օ��������/�+Q�Z۱tAO��F6�56�t��I^%�\�Iڃ%y���D��h*i���}�.�e����PSC���:���=dz Q6����*� tK���s>���HR���@M��N;��c`%j:�c���Xnƈ�>����#��z--�I��� �;��*b��2�'�#�R$��-����������x�]�
�1��+��>[��m>�-�߮�9p����h�-�ڭ��,�FW���d྄�&���i�P�b���(�����̻P��7$)6��>c�� ��@=�e��U���� v���,|��ݴ��5��x�šP��[���aK���
��!��^���c�>Jb��CK�
шߔ���H��î7��bM��� ]���ͤR���w��V��s�����:�������+�_/����-���� ����"��=�-d�A���P1��~���Gl�7���6�xg����/�`A���H����ɱ��ފE�H� A�=m�ݰ��Rp�&�UcS_�8���nЖ�n9��au�m�!�k .^�����_J���QVUN�1
.<vh7�o���Es�WYѥ��@y,� �a�E�'9`$)�O[ʀ��ή�[�@O��=�U����^`Ą�8T�uЕ��|uO��ؚk5�k9���V^^TL*'e#��a�5���Apǿ	�Oa��������5!^ޤ��">���t�t�pxo�A��3nV@ՠw�FF�x�%��;�u����Of���11����������2�7�GQ�d�G�C��U������+T��|�+/^����XZX@G/�N�6���	�.�z,'���:��EJ�7����$�z,��BC�A8<?���K3pH�9O�Ș��#	 �T�����Pۼ�VU`֘n��SeR<��ص좏zL�����������2���daz:�21@2Y��a�. pF���ƝsG��&�z߄��<NKC-����?k�^^M���M`J8�<��C_�M}?Z���+D:7�!�<����)ͱ�|C)�G\� Q�ߨa5^m���=M6� 2�c���rr��K	�_�{���;Y[�)ݶt�fYZ����gC	@'[9;4�4�� C�xyy�d�ͅ�Y������j��&B�r�:�%}�A�)��bG���R��/]RR����cL�jgg7�e~cֹ�J"v��J�Jچ�߼��V'H	�Ywi &G
�����'���e���y-���0(��wa�4�%���q��/4�8x��(HlO��7��#P�����s܋H��y��&���b�k�T�{%e�ӵ��M�sw�&��,��Ӕr��ąn]$ ,��ĵ}������R�ٳg�L+��п=F��-����n(@u�������d���]�ѸE�⩇��=�>���2@�Th�x�� ��:I��RF��,�X;���2�n;Pr%���.��wQ�.ll���J#j��)����y
,T��R:�?^��/�4 q s=@����%(Xbs��E"?���V��9Z�Fu�����Y�3��9�ctK/G!(���3��he�𒖖���#��׻tt^��ns���]Vb��T����KD,���ܪnn��C%��J7,��~��I�������2��ƿFio�X�V��oK�L�l&y�����C���g&��xy݇vD������i�l�A�&Z�2~,���� ����P����񳖺�^bku+���_9�VP�|$�-m����>��M�ޯ5㸍�f	��䏛�nF�}�)/@ό�E���$$$�VV�6�4��ٵuff����m��P��m=;;�r��1��,���ЧC)������Ȥ�� C�]�������Jo������&{2��Vxxx�)=,/��8%�IO����k�ptMeL}��f�gK�?Sq#���4�������§y%�hN66����ԣ�>O�꠴��ܳ�ć��s���g�`�lo�܌�pu�����s�<Z�-�V̇P��`��|����weeZ�i��q��g�^���B-S�,L��3i�_����#N\Pb�˖����	(��8��_~����*�,c�6)J���p��� �1�y�gg��3�ffߝ~��������؜:�������22XI�?y��j���ۍ���ө wX=�3�'`�GS�*��!	`���#��&�B��c���)�Ig�N�?(|��|�U&��,�} ��)���w�@߁b��@�X_[JᲒ�����?�*��h���9:��{�uq+�{r���>Q����BzE��������^���\U��@_�����n������{�M���y5j��8�+P�Q������@� �<��g�d1x$P�$���=xP0(��)�B_����VQ*���&
��榚��{]ݱ��Қ��ax��w�;G��"��^hm�ƫ��4u���y8=.�,m,�2_�������*���[Q��w�\��P�����VNBD���� �2Kn��]��_��U��>�F����6�E��p��i�e�EJX���|aikz����Ďì�{2ǃ��W��O�kk�����^�)(( ^Vur�|Q�P����� r��4��7cv��]�4E�?��&h�aL쥏�^3ζ�!�ݛ�m=\���Pu�qY����xJ �*�<V�N��E����HEق��f��$�{��\q+!_����*�*�����(�Rr��g�zJ�#��#�$$͋�:	��K�T�O-hN�9�nn�&^SEw#�ofdy	���
��ڝz�t��nL>X�O�E�i���6S�~���1�i��Nrڨ˹E&Ũ�_� ߀K�j�����a�<��_�6y�[bE-�!��K���*-9򂂗�B�{�τ@�����uK����\27�߷���:�2��PHH�6���S��־����G�������P�=K8���7)�����O�^Q[�ݟpI���k$HЬ�ڲ4��F�8Y>M�A���Q3��K�à���6����K���� ���%�� ����g-{����'��)��-X��3��)�W��߽>9��^�Oo����މM���z��q+<K0�9��7����3�^ٍp�0w�*���{F.��ι������ﾃ��� �/�d�c
h'ܐ̵�����s�S`��5��twx~����0M��c����!he^Fu��P.��G�ed�.� �o��r��Pu(eV$��g���4˵�ʵ�">W0A�cxxg��Qu�_��0sr���;��L�E&�b�?5IFD�-��]x��"rI�e�L�����겇���!�\�T7���HNo��o'�b>�APD��x�'������C
��w����O2M0���O�����b�2��Xߵ� ��F ��� ˈ^�퇍���LR&�[)h"c�p�l�:��5����K��ؗ$^���R�׬4`vh�� �z)"cpZ�{�T�\˺3l���
�(��X,B��o7p���7E,ۀd�e�Gl�X�M�Đ�A\nB��a�d���4����I{S�`C��]���(&kJ�y��-��Jk�����,DQ���Z�--��w���h��H���,Ӄ Rl�ЂG��6�³ #����Ng��axI��Z���N3�n����#	��F�8b����\�p���E:(o.*V��L��t��G�
}��zG���i )�A�W7=�r�0h�H�k`�x�噥"YO_�[ )d�۔n�(��S9"�ɁLhY�fYM���9��<jʔ�>g��/��˦>��'�U�K�d�S�\�8�ʰ~.-%�D���!���\=���[ )���
�����^��>�����v�?�tz��8j�Yv�id4��*oʃ���?����s�[���2xJ�/�P*�����θy�͌�]X���������;ؒ��6%jŘ�p׵Z��|�:�9���=h��'o���������κE�l������TU6.f����^щr=�ˋx�&I	�y	x�fR8/J��{�k�5��Jì�C�#��IVƔ���w��%�bc��
y�K�fӂ��I�[��ٓ�+ʌ�dnQ0��T���� ~n]��y͸f�]b�F��nuuI�e�8K͸>6#��]~jc*���c��92l����﹎w���I��&�ȯ�����n��,�E1��k{F�))� A���K?��,�PJ>��.��Q�����&@U;9��y`������1�gx.�[���ǺR���-]qz���ԁ��ԙ�欪�P��C�N�L�]���]
B޴qAte�T�XҺ��c�CN�t�&����Ƶ0����:������g���ɂ���8�E����T�j�*=�u;�R+9$$HΕ@0��+�HH�IB���Թ֚����@�c�/2�_}O�^�s:${���h(^Bۇ����||N���� �Y�ԯ��Ȝ�I�;��_�%w7잒�}�z8�?�'DE�+_,+j��2%��Q�s���Z�j��-�C�:&��ȱ��.��5J-�in��ʢ�)�'�w����P�X��R�	�}zd�Uզ�5>���+�Vѻ�c�x��;e�˼Lr�G%�,�Aᳬ�ni-���������j珘n����=1>D�{R%�4f�1�5��K�ϳj�v��|RE��Û�lB�tsS�y����j�����W.���/6��cN���Y�GK�E�;f�i�/#B6]����n������v��Q	�ѿ}�"��l}��6��A�P��H��ZJs��H�V_���l$^-��?��X��W��t�|w@�75�nFV��ωԛg|�j�`@Q$��%,&=$l$t�����S�(��u�`4]d�&�'d�G�o����q�?>�
��_TSx��g��:��=�mRp1����^D�U*����_�ñ�oM}����ΆQ6��2�����}� C0�+o�r�}NG��4m=}ve�^R����w�w�v��o}�����i����Y�X�MJ�Y;1P8��EJ���c�jsN�5���eNB�ߌm0|+�ۻ$������8�͓�?�N׻��\� �L�;��0�c���,��(�S��p|�ʜ���5`{DR��2��kԜsвZ�!~p͙t���N����'M���-'?��jrz\���D��6�����Q�����%>�]~nl$ZMM���ڹ�Th��1���p%	"�V=V���=
�,��e��0?����_~ԗ+lp�ʴ�O�O:%���Йoz�C������g��HG��)f?OuĦ4-�X63"�$� h�?!]���^�HM�FQ�m��׈e����/,`��D���KHJR��J�`�	@�]ZR��o����xz����������IvV�i��D�[����s��m�{ٴh��\!ݺ袹s�Cn��Um�sL�����+ � .//_!e�!@��&8�Ü3]w�C�ϣ43��H ����N�KHD���^ZZ�r�e���|��Q�oT���(ŅWI��kX,a&T,���&�W>�9�~�V�|�-�=44.nm�4??���rWBJ�9���5?h˴���֖���(�k��DDD��u�&�𖉡��T���*Nܟ���N�\1�<I����"����q-�r�N��p��5�;�ql2J�[O���UU�����~� 9P�%Y)g�\H�too���D��o����Nd\\\�<��B��;R�t͡�u����}�~I���z�KP|씠d(�aƚ���#$*̒�v��C^%�޴�V�q�]���9CwaI<���Q�W�X��eV77%@l����w����t�����#��8ݟ���L� �o�K^��|I	��m���6"s�>��.!�M����fRhh��R��(���x�Q��;�?n{�����p �Zfyl|<;/�N||��u����j��"�/z�*��}�)��ەr�Ya;�!JF����Y�1�Z�]��iM|�p[T�ٙ3&&�]zz$*>9;�#n�G�A��������������Ȋ
���Ĝ�\��].�^�웟.���Tb5^�a�B˥��F����{��|�Pי��ꇉ�
ntj��P�G�TT�`� KX�ß{xxd�Y"�>I��,��M}ਯ�oEHGG�+��72P�F��(F�.�/3���QZ�aqͲ������J�wd��ۜ�R|�V>���wycccr

�����%��)s�+M��ss�@��>�W~�Q;�E��H�.�e3������r�:�q��ylE�ō#ﰣ3>�A��D��*N�4���{ڄ:�ث�U�RR�===`>��r`ή���{<Zi̙���ܛ��EFb�
�����&=س>�����Tޟ�a��U�`&h�Xr6LI"*�y����Z�s�]���F���Opg�UL��C+�?�N��:��+|�q��$�"alL�<�u�"s?��{Cè��;���hWa��C�����>6���ڊ]��(w}�8��du�7�fV�O|Jg!g���qtt|����iF��Q�:,4TT^�t �I����^���M1] tyyY����Vl�S){���QRl�h��b|iz��Y�t��d�C|���1u�.=9[�Q��{���8,|���}�\4F�")!�|g�9I���)r\w����1����z
ۇr�V)�451-(N�Ho��e�kb%��K���DO�-Ĝ�xLz��׈���SE�����&����5F��j�u=������`"	&���9�f���rr����3��M��M�<��e��o~��>�� ���~�E�w�	s������+vVY��KN~��_���wqᵸ���:��;���q񮬬,��0R���C�|� >�y��r9; |7�Vo��$S$I�LPK�T�5�k-�� v��!���9@/��1�x.HsKK�g��M��jk����,,�2����3̼x�)����ɘ��d��N���m/�,����@�a���rww��Z��R���ۏ���g|�~�6���H�b����� �����[���8|�χq�J�|���S�s	<=����T�Y�dR�((���[ɥ�n��fgf�F򕤍�?<xv'1)��ɰ��7�����
6
*����C�J|���ũ`�k��W1-G�Qz!Yśaˡ�����Ŋ���K�̽���U�g>�������S��Z��_2���m�@�k���	cv��
��Ǡn+�����,.��?����>�mT9����2<İ=��;ra�jkr�wH�DK���ˀ�(���or<6�'^\\ɺ{U��4�Mz:)(ٞK'|i��
�?�����?;XM�id<�3����~����~k;�s�Se��λ���`t44H��$��$;;�)��H!&�\�DI++F(<ZZ!�|���&��{���M���{�bI���~�f�vv�j;�T��G���5�_�C�n]��to���$�l���_⣐��V��1�Z�Wg�����G��ض��U*o���
�����oj�Ѕ.�m�k1g�M�ؖ\hT"w�<ƪ�xr�!"J'B�,{y�8�q>\t�l�Kh������1����Hb��j�s�±u�9�bFe=��55���T�$�W&��e3S�{r�5��a+�����N	>@T�t�Stl�B�s3�h�z��X�﫩��Q�42��t�l=��t�^t��k��I��p�,����}�G_)��(b(�Ia�����+�+�iʞf5�&�� ���+ʅ�?Q�v��سS>>&k��|�~�M�Bmmm�P<�Vv���H�we��L'��~���s�W܊B�?�S�"
|�l�İ4���Ո(x�$���e�aw;m훰��������h̚��'���EH�����>ɗ/�"Ʉ#����\v
��KW��:BR�g�CC����F//��/P�1KOcb��z_�k��)�q���R03�k�9 m����ݲ�˯W.*���3� ��B�+�z4/`C^����}� Gh��Ej����ݓ�i�?,x�����)���D"���£�?B�Ȉ�H)����e)P��|�w�d���J��i�GB�����D���4:&&�Ouk�#saA�d��y]ؼ���(�5A��-W�����宮���p֯��Nb-��zz�� _�]]T@Q:��w��>r�8q�a]�r<�&�������P����`��+)���p��� �4'
o�������r�SG���
ç�|$	,�a4r	�uu�n�_@��8޷�iL3�=%�:j
{S='��N��PHQA�@���6���?i��������'�~��D����~K�fR�ؓ�%&C� K��\�h`���P�l�ԛ����b���P�or�G���	�̬�y�H��U���s�+!�gӾS7�9�J~n����%:::?�0�����܁h��t����G(O�}���hr4���N�q�N+����u9
r�N3���kp^l��^o`?���.K�Uc`s��+֩FED���k�ۀ-�=B{��|l���O�6p�PB+�	���I���=�GEy��<b��x��T��$��^� �!v�Y��iA�ѫCQN�]�n�	?�����6S��I��Y�-�������;ý}�E��Ǳ*��c5Q�Y�߸ێL�V'� =����5�"���`>���Ob�9]��\>�,*Z�ɗO��cm�]�:�kSQW�S^:��Sc�~�>`*�Çے�����G�	��9{�z��Y�BM�Dw��9t=��s�_�!"C��a?�i��D���ZB�k�i���R�}�m�����J�Ԅ��5��[���$0����~G\�e8���0�(1��R�0��쑉K��> n(f��}�=g����CC������-�r��������;,̍Đ"1���?�r�)_�r젓�����~m�׋�Ť�e�	�1H����~�òCRS��S8�uE�u� �{7�m��oT�\I�;!F�Y>�aV��ĝ��`���问�Ej���5{h�b��5��%%�0��@G��(���{}���S:��'~�͎b-,��UL��}�Y��_���n�����?̼��J�!~�!
��DV(�л��\�;|���"��(�����nZZ��i���H�YzYʐ�z�*��'NBt �?�Q���n:�}c�_��~��ƌ9��޾�Ty����Q�y��=��<�o�]�
xhP�O�oC=tϗ�~N����/.�CBC�T>����~߷�X�L$��"zNNN�Q�,N8:B���|o�X_��ج:Ռ�U�^�tP��Jďϱ݊�t��K�R�
������	�ne���x	��R�үY����2Z�lht����� �ɽ�
AHC���*�(0Y+Jo�!u2�0>�_J�a<(�͛5,�	%���.���;ctg>$A�'��UnZ^齆1iOt���Asp��K��q,�`�����T�m�{}j�)̜`L�f���-�=n��n7�.���j�֏��*�����9��
�YrA� ��֣�}��}�����]�8?����c�/��%O��#;�1��k�gt?!�`�EP�k�g$��f$9���h����'S-A�N˷�ẑ����Q���r��3K&''O.�T���ܳ�r�W�V���w?��&��k;H��67������M�Л�o�wo�t�p�NV����i�{NL�`�S�D�fa�s���k���^�,'��v���M��uT��HJ��L��ۙv	�P��𯫜����n!��Bmj$pB�O��鲛�����^��� �UwyWQU���sqq!]�o�;���A���ХCR��%0�Eu�>�^�;�6��HS�H�7���S�e|r�����s� �
JK�n�4���5��������z�����=�o;�,�*C���+��'���>�@�y�E6ѳ�b������^�o�i�{���-YW�˼9{6,��բ���4n�<�	����a�w�P^ٜH���v���w	-spq���g��Rt����x.
����bï�������H�Z��S�f��gcHoƘ�?GNM���r�>!Y�R���]{�.�������d�Q��ɀ����U+��u���oAÔ����1s[�ga�p��;��?)3���(X#�E�Xb�52��r��'T���T*6����v�#ԼΣw+^T�ߑ�o��N)��Y:��r|D�����*䴟�(}4l@����p�$����Y�Le:�$�ņ��_�<�E�$4�t�(���0���X����*ue��K����R���#���W$�V��<����tku������x�-�^H����Cl�\+W�h�ɝ@�G�uk*h���;x��=U��z��+,���-#g���\�J��{{zځ����Y�1^�u�n�+Q��/���߽斖�y�l�6VKOn-�6�}�s�J�	�7�M�����k�wK����Iv+"�������=t���-7at���d�%W�]TԎ����c�_���m̵��ב�o���օy>۽-�[z���֩i�z}\IH�`
���n����#�α5Q��`=�n;X�8�Ǳ���|/,����s���A�r�	ޠ|Z�W�j�1~�!��f�M�vC��5к@��[�1�d���O�WZX�|�����;52�_wH���CS�o�S�5 ����|a!��Hr�w�>�
���u䷕4-�v0l�\���~sNª��O\򧧧I��<����:��8knw��H-o��S��G��wO,i�m"<�>�s�/#+�y��}tz�v�s�/K��{�񲸸���� a�f��lc��ϵ�|���cy��q�F@L�J+��!�(��>����B��P�S���`�̬����%�C9����Ƴg�pϞ
S�d?��u쎇�5�6R�����*������� /qpۍ�- �Xئc�Y��A��e�JјV�+6v��\P��1j����`bv)pϼy�a�s)��Hk�Y{J��R.�k	3�n�`������f�zL�x|\'���&�\� �f�ߠ��-�)�N��A�~�kVC����'I�o.���Ѝ���79E���Lq�ǁ 7�ֱ����_86bGQ�����|o��
��u�w��B����9��JF�����8	\�oD����
Z�F�f｟Y�!���a�L{���e�7�,?HX|����}�B"o��*뢐�Hhϡ���˗`ʃ��Shc�uvvv����e&ddD�}�&p}�O�̼��"g-�h};"߯I��>����!238}B8w���$O�c[��q=�=�Q�2�tJ(��Mȁ�H���V�Һ��1�XDh	@�ORv�?�`"	*�e���+���-�G����#��
�E7X�Ơ���-}x�I:��&�����	^� �ң���]Lȭ48s�L�ߊ@H��p��= �\1��sQ�	��V)�/Q�U�i����BDW���.T�]6�EW��"��~#��4/����k�wy��wZL@�hs<''�u��n-C�20 /����}X�q��)��bf���>*`�r��9s-��_8K�]x��Y}�Y<((�d^X�ؑv���6`��]���4�sK�uZ�L���9��u0�@�EAJ`��w�_�?.�1�����*��[:�s-$R9C��)<{?��5Iw�H~9�Ld�t���u9���܎n����VR�R>Pz�һEo���s_��^wSt�|��pͤU�y����.$2.rrWy4Z��� ������ZQ?��������d��[�v�U��w~Y��ꞷ�ͽo,�f�?ź��'x�����?j���(Qq��bO�G�$��j���3M��yw�~���i-������)�(��,h9�E|�L?���P��zd O�*~��齅�K�.�F8��8t��e�PX'����d�T�)�����gi>�v�/��C��jU[���Π�)�8(�g'����))J��%L��K�
ls>�e�{��4Ү���r��;_:;Oy��W=6�slba=Ɵ��N�W<��@A D3t0T���|�/�%*��9n��C+��}<���uΣm_TX���Ə"��E/��l������C���g��B{l�WύZ�ba����� T]��C����48��Α�eϲ�"wsG1c2�t�?���J�K���Ç�3.��B+�FFFEE�no�e�o
�k�ó�邳KhK��4�'�<*G'&���HV�:,~�M	�7Q�H���	z��}}�ax��j���,���
�-��؇e6;V<�ݖu%$�]�*_�Љ�/'�ϫ8�����g=�W�g�B��X%�fd�Q� 
��������V��k�s�@�k5{p�ZVc�"a䪆��<�z�����HX���д<p|��D��U���_�[�q���=?�
�6JĲv�~�����1�m�� ��\-`�^n]{����z먪��_���8t�N��D���;�	E��� ���%�������{���d8{�91�\k�H��d�6SR�;'ȅ��P�5?���/"�t�+��eRg��]o�g:��Qi���;d((��R}�c՞gf�s��/��F��ӷvv6W�c������ζ�nj��	�]�i��h(�xS�'�	�����z<���"f���rbb�q��㢌���t�A�M)}}��"cc�S����6-��#"m*[�)��/oz,�e Qc"~�O����h�^���Dn"��+ �O<T���100|3X�������
�^���x����EYpa����Rr�l�\A��<���l��j���a,�(�"�t��ܟn�$4,��Ċ**G�0�腋�dߊ�����at�ׯ_�r�᎑{(����a��i+e���ݍwFB�V����]�w��8� ��EԋU^���n�� ���a�O^�qb8u]�����\���'�N�+v�H��mfL|�����n�;s0aO���Z�D;c�k�����d���'��q�j������r�8w�%/���r����P�J1����g߿��O��z�Ժ��'vc�w�@7�qǭu��ohh�a����	����������PI��t��%�������]ZIC?�MQ�9Q�|�}#<����>j������q���� �_n_O�iVW��:�?ߗ%���$\r���|���$%�)��/r��)�`�w��#4�ū,�~��@�)k# �����wm<�hN��y۩���so���䎌�J|h��z_�xq�|�O����H,
x�W�J�����סEC�_���jk\mr���ui�����W�}�.�Հ,dL7@����-z�@hA=������_��_^�,ں��o~0nxF����;���+Qh))�Z'i,^W\ ��R.Z��ԕ%�|"a�KD�� ����I�r��/0Ub�p`&�s�/үa�����U�ݨ�`�h�~��=$id��K��X 8c)�FW5���;�:��T+lll���ݎh��oF�p&#J�)�unl�y;����!.N�����2�q��=WQ �Y9�1��P$O��U���
�������zw���;�ߜ���<�X���� /l��#'ߥF'�j3d��+r����@�J;;;�c.D�+}��Z�Ϝ� ��'��<��,�[J�K4����S����6$څB���r�����y�9��Cw��y��*wQ���4.phZ�}��4��|�j�o�,|�9_h�0Z��fМ0Z5��-��9O�.��M��}P�*��RS��ø�5;����X�>���$�nc��+�~w�4LF��o�B�=�4˦a���!�%�٢�iNwB2�1���(�H�-Y�'�\���r���`��/19����Du�K����.r�?8�Cb(�<ɶ +	 ���p��u��X�W��ͧhK����������|���-)>~PE��i'j��ye��������u��m��|1u��;������i)�׈/�}�x��6���6��Y덏���������*�P��QI{;�L&=��0�ri3��T~42Z��^KIn��.M��/e��9=j�*�C4���ɝ�X���ӵ��f��8��}=�7���2D\��lm/-Q��F� ����߾�HH!��5'e�R���Ӻ�^ڢ��y�kg���rsss]{9� vi�|����-HJx��#t�R��(ȱR���+��KGo����~�ohV�d}�9ө����IJP��llN�[�aS������jj��;�a��:C���عM.l%.R3?���>�u�Y�h .=l���8O��e�Y(&��5�g�~��	%�U����,�o���IͶ�kE�Ԓ�� o�^��"��`0�X'!��[�П,x�*�id����2���܅p��G���ߨJ��!�p�[�hO��}.jv��Ƈ,n;��#<+��f2;1_2�����	�N�pb��(L������}Y�m�f? 1��V��1�n),�w�WH&�98�1��L
�A55�c:/������^��;> �����<v��@�ߗ5{��1�؁�|Ř$jQ�ޠ�D�G��!����3)��
��lQq*Q���G��h�;{��d:�̈�3���3��s5V��z�(��*�TTS�;jX�/�������L�Y�[px6Ľ>��Ո_�A��d�JBW'�@�_�������D����]vE�ϾO�A`�P���������	���a��d��MŴ��*P�yQ��|��)���Eڧs�P�m�K��}�M���n�B��(LL�
����~G(A�3u�F��NN��?=u<��A�!�|s"	1qx�IE��HOOo���]0������>7�ٲ���Ѯuu���*/j���k�Ȯm5Cd}�׹<٪v��tLL��ғ�gֱ�)����T���TWPZZ:�ĺ(�\�:$W�����)#����A�{���:�_�(��)[�#Z����Omzz{�s�*0��9~�� $HW(:AbN���9�3�Ъ/��ぱ�����0�x����\�H��.��b֑[�%�h��*��/��W
aHt�p����5�> �L̛�����Gǹ.QuW��<Q���պ�O$V����q��n��]�JG���ŗ���"��T��A���BF�7����ҡ�"�HOn�\�j	D)�i~�0ڰ��r���9��w��[��t��/V�fN's���Z�zO#?�U���g%���N���� ��
Q��KCӯ��Zw��������S���K�^yo��J�Ԕ��7��"#מ�t&[��!�+�����_[��Tr�r0����0�Z�Q��g����S��0h��0{R��`�����۷�r$R�E4o2��`�F--����-�(q��'K`�2��a���v�n�җ�P%wO������EO�� �zG�lv�;��d��/�x.V���-��Z���RY�p�ka�BT:���KZ��� F�<�%Rs��U�Ȼ���F["Bm�����|���Pv�;� fL�`�NBd^B���Ng�h��ѥ���	qT�¿�
�����p%d*~��W�e�X����ETT���z#�2��y�¶D=Ry:M�i������ܗj�Ҥ�/i��bTf-NO#�� [,�\?��������\�B�4G-���ѐ� ��O#�K�����̃����ZWY�9`� ����e#���A싧
��=�w�ݪ�7�;8��6�a;t�$K�%u)���lؖ�Y4����ǿ)�s�̓�E��[�sttt�qL�x� B��+'���.��S����'f��#s���g�YL�
'q{{ۯ���a(�5��H�Vm犺�q��n�|��^�����rH�b�z��l�u ����,��$e͵��~�]��m}���|���ɇ��x�	䰄ҳ��3t�nn�pm:�6v(P�
�І3�[7���Y�o|�e�����P�+N�� g��A��*�Vu(�b�A��hBZq(����}EH"o�G:tG>m���j��6�� ����I�����w�I %niJ���=f�t4��
d���$$!���d5�GA�n��"�Һ��M/FG��/�V�D7���:�4Ti�VP��^GwW6����F��"��+�c<lU@^�2���%��\�?�gY�4t�qeєg���=���c#@;��沐Ϗu�B�N��Pq�ũ��]�0�3���AߵX�ߗ��[GGU_�<e�������0��`���ޫ.ّ&����ַ)CP|�罴��XF�1�2d�Ǐ���T���,�L��jg<2��)�I%|Æ"�����!$����H��F�H�[��mXf+�h�b�s:�%����x��1@�N���(<8�۾�������U��0@��A�Z�:���
�q�I=�繁�����'��U;��u�)��������<~s�000�ؼ���;�u�����Z����w�ҺX&�YwVu!P}�2kl^��ɕ��6p
�yV��e{��8R��0�v3�
���d�͏��F�ER�Py�R�to6q�8��{��L��;��Yב��ʊ�����*<��~6���5���+�Z��Ax� @��Fv���\\�
	�G.=�!jx5{�h��jLC��S����$[]�����Z~���8����;���ިYe�)���e2�fA@}�Y���3,�_�ˁ �G�V�O:��r�o�v���ػc�fP��X��D�h�6���E�ѯ�tL�E�4S���7�8�E�F*��K��q/�����3J�T��8��H0�Fbe���FvbL���o�����߾�J�����Ǆ�_x�O�t�|(?\0����\N��l�+�tc|;��Zf�,~�΅���zn�cs����8$����/��v�h�X����H��"���9��f| ��8K��.�u�*�K�g�PV������Fb`�}!�a�fKvtry��F	���l���144��di{$�TK}�2�'��=����B��0���6,p�g>��KGk�f`�R'u�X-��x�>}�*H)��~��!�w7i�����O?����=k*�0�� ��d87���h<�܆F@�6+�up�R�v��0�‎:�	�m��o'��f8�qF	��l_y4>�꽂�t���o�F�Uqa�U6#3<����UGͅ�ƿ��������p�)����Փezz��o�c��~����N�OI^�!8��8ݜ������F47c'MrQ��W�{�_�`,9qg���g���V��Q:w1N������W#0�FFF��m����3��F#�G9��*
 ъհ�uXay�L�Y��s���$S����n�dz��O�aSl��	�}�m7f/���' �,�����w�TY����Ĵ�p��k���	�i��LR��n:}i��s�o�D�d�*�{R�c��O֖蚶��M��Q�͎��D���� $�g)G�~�������{�B��o�~��W��Zl3#q$�Ja24�0�Aa�!R�c�<"���S �*�P-��C��Y��b�V�J%����%�Gb�I���S���/�){#jI����}(3l�+���bR301�����;WOV�NJMOg``�^���r����p����C�я�j᜖�y	���UBi����L�W���qs����3)��M�A�s�v��J��� �-��EN}�*��`e�g~�ޣ�Tz^�i&߃k
�;N��޸���O�<cbwOz��i=��$��|�VU�O �*~�=��wǿS,s���{{��/��32HA��$$P2>�g4�� ^ۏ�e�p&?���O����}�nD�2��3B_e��o5�|��X����O=����jg��T'8�t��Kdx���HM���7`�0a��v��7QE;,!�q�هD��dD>T$P�ľD��L�y����m[-��T=6�됿ӛ��_ZQ$9��F�^���NF{a,J��Ą��I.�E5.~�	��&r_��s&{-�4���2|2t=ɖ8��3�Aڌ�9�����@2�5���8��;��_��<�+q?��!)�E�b����藄��=�Y�|���fJؒ.O�@$!X�/�"��vajBT[SUB�<�Ǌ�b�$��2?���Ʌ�U)��X���ܤ-np*Lʒvv���͆��,�!=��S]������.��|�GsVzR�m��3ާq�τ� h�����K[bѩZ�n��f e���!���aB"��Û�x�6R�
��C?��S�]���GW������j�A�$�4֮���jEA��#�F�JW_Q�YyR���9߬�4,D���V�v=M�>�=��|j��ebzZ�+~! �d"pn����ꁷ�Цe���FM�v�/=a�y1QmE��Yxxq漿a`����/|ն�/�) ���%�J����w����:�޽`c� e�r��HV���h�0����4f�_��G���1����0j�{;0%&&�/#���d�x��E�C���S��I}C�����}�#YD�����u��*� V�������i�7�q���-]S���!j�"J�
%��w}P_��<���w|]n��S�q�lB�|y�6�9��$	��7
`Et�!;Z���s:�5;b�Z�:��Q�D�����ӟ���<͓�*a���c��g�������(�h�Li��V�5�w��W��C���$�Vp�C���΄�Z����bc�N��/cj���F%C�	x�|����Y���!n?�)�+w��޸���<���42	l�J�l�AQT��k��0��ܘ�.a ���% �x������M�w�=�#�~ư���k��ڪ|���ƽ[؍qJ���� �O1Lc�T3+�K�u�ؗ:�N]��cD�umC���Xԫ��=C�\A�MD��A�_qЖRD�В�"kv���G���>>��ĩ���%�ޅX���O}�Q� �� 	�i2�n},��:di"�#Vu��dĘ'e���(1����M՜WdGGK��/?�ج�C�19����C2�����m���e	^�n5�>�x�#�$��/��wi�E��0���󋘃��?yl[�dR�[Y%����$����k.ܼ���MC�$0A\;��S�L�t��ưi[)s��M���HWPP�����U�
����KQ@�܂q�� ��l{�}:�k�"��` �����g#�@�ȑ�[]�Sԫu�c�����Œ��>&��}R��'RW)��Y5���b�]�	��C���JV?����"n,��j7��=�\5$1��Dv�&�I^K���M2F��Wv_и]"�	���2SЎ|����Ew�֜���қ�g�$�Ӹ�m�(���s{��R�ECb�/3�x�J�$F���J�����uH�u��|����j���\d��A���Y�r����8Z���J������v-�_��Rh�NPѼͤX�\���ݜm���c)3���c��;���������.ڹ��>揄>�&]٪d���FIuEm|�tL���>j��b�Ng�5��yK޸Z�#f����{���4�(1:�%���8�_����=�5���I;m
��'�P�HڋkZ�v-\�u�!4""a���Uz���:��M��#��~v���J���.6�KKt �C�\�b�H?��Ks#j�(�I�Յ��RNFF����-�Ĝ�Z�q����2�߫ݨ��Wͤ;4�+�������V��~>h7��k�Ң��r�J*6�I���1�Sn��S1�������~+�.Bm��M����S�uJ��׶�N��;����#~�.n�<������~;=��<�x��������n��.��l��c�;���y��HO/Z��UK���/J��oY����i���%�w=���7��cT������{�2�bs��]��E�Έ����@��9]�?z{��@��r����N�OŮ=�9ۂ�>��^'�uB���u^�q������Ԏ+�� �.8�*�$��o�$V���8��ʯ�NO�:�+k�hR�lB�!��~5���=7���w^�
���Qu�×^�;����e`���^`{i��%3l�n���'&�(q�am�A��6k�V$ ��8 %wn;�V�̳�����}|���Z
@�G���u�����ป�_e��x��� ��Z���t��곯�W ^X�|L��P8 0�ǫ�̙8[>_���.��Lj����ȥ�d�@=οa61OH�R��_����r��kbIK�J��;�����/����w�d`o�l"B�[qg~X��Ki.�����0@��o^8<ɫu돗���$>-�g�!LRDjXvϴ+�@	o���FI	�i�y^����xnf>7����t���V�����4z��R:[����D���6X?�!���r�ʢ/�
�ƖB�P�������vY���vP�M���9�������:����h���Q;��|�OO<�sx�dm�	�Ɨ�F�_��t�\�*>��34C�H3�w/ց���o����#�A,�]v�[���#_Y8��-qb���=>��CG�QrJ���м����{���87�w'�+NBxh��2^���l�=E�bO2�'�B�)S��un�(̽e���;��;�*�yZ�}�ϥ#Ę�n��

��O�g��cc;�8��;���Z������|��u�=N�&b��{sZ���6������Iol����Q-E%%
�-f�(�	=��Rz������|���f��=rg'E%F�~/����U��k(�ۑ�����.�&��)���9��<<��W�Y� %��8́��F�<!��%�=z�����F'S�%Jp'��K/�8�KJI��$�0��d?��*���>��S��1���s:�[���A���}��/�w��DE2�*#��Z�2���ʱ��֨�^s���[������Bl�ջ2{�	���%��l�uǂ�%���n:(�tD��������C�w%�N�z��(�ꩩ�jU���`���:p���l�|�=E�~����P�U�\�)9��Y������g0�Q�LNV�q�����W]��J��?'���ݴsS������gf��� ���y��eg�s!��/8�.����꒴6m����������Ӡ<�-�.<�p�	�;����մ6%�ڶ8Rp'm<�X���u^EŨ�$a����a�G�&U�|�C�7�2�/���x�M\�U�����é�4�Rl�On�IX,;q,�zBo,[ք̵�z�?��/��u�҈��������ޠ��^ ����%�ǒ��G���$�|�'�S�l+� �Ó9h~-���sR�?@���,�l�Mx���T2L{��Rc�9�Qy��x]��WV�Uo�H���B���hhi�2*��Z�ir;�!=sGz��RJg�.�O���;�W��l�	����y��=t(>��È�3�»w�&��BB�W����/yoc\��}��r����G��b�������N���S�P�>Z��˧�46N�?i�IR�}�R�`��Fr�6�to",�8\����?��纐=3�k���y}��*$䵗����#�Ǔ'�5�d����8���W��)ݥ���ѼSJ��aGx��Ir,ED;�����I���C��7�X�����W��.Bˮ����b����T/d��rp���t�;U|\_/���� ;A��cc`��GeR.A�ov��d�y�)vH�Fiz׽DK�D����L���i�pi:�q�ϟ?�J���yOV������2�E��T(CP�7�Z���Ozj�������Q�
 ������=M��Sݝ2Yy��]���j,�Ǐ��>�>�w�{��L�^N�nk�F.9B��= ؘ���↘�|ܶ�k��F��u'�k�V�[��f�'�$m\(��`�m<�%t���B�{03�_U&�8.��h�A�� Y�ˀv81�z�<�(���}cƺ�QZ����֤���T�yӳ��J�Td���gxcdw"VXNN��ǟ��b/�?��R{��O�ёǽQ�‍���Q� 	T�T���;(r�c���� ?Y0[.T��%��1�t��e��Hz:��QC�_��ͳ���0�wZZk�I:5���o�T�XYX`�����U���߫�t��%�GMe�Wl9^�|�5���!�����Ru7m2�)�&ks���+�Q�<t�����6�(7d�A��1�����+t�ur��m
��W;�����|�{���� ����_f�wn�}�!��/(@ڨd
�k$��()aifw{X���V� �av��xh�%m���P<����`�B�l���<���>���kk��z[�M�x��{n/8N��\\j�[�p����rb`����R7o���'|]�.X�m�nШ.]�TdMN��Vo���u�O�g>��/����4e/����q�e�_�n�|�o��R����'�Z�K�͚�򌠂�	�p4�����_��,�K ��$H���e�V��k���!����	)LԾ�U?i�hC��MU�y�
4�bׅ qppTl�L��S��.��#���Q
�_Y_+t54x�+����������5h�PHa�9�9i�󺻀��`Q6��ဖ@",���_ c7j!uss�zt��h��@"bϚ��Ӏ�N�����v�$|����O��vs2����̚�fC6C�:��\x<���s���|p�ͤ��F\LDfu2���"��P�]zHW2X�(��_I6Aw���p��ap�
�v4�|MO\'u�]H��~q6)�Ŋ!ٺ�9N}�B���O���"_)�A�n�B�.�肵}715�ݽ�h&��F��,�<���� ��9Jlr��|h�I �;n��Ov��?5�d��'� ~�DAE��M�$� '������E����� q���"H�T��c����͗o^�*��Pq��[�Io7���Up6'%���')l8'�fWSCEC6񾰰��P\�4������x���yCw𥚎}(�3��1�.�����m��I��cq�	�g��D�H�o�om�3��e��#�T���M��*��B�N4��ݯb%.��[�^WU�AH� 6C���`gi��	�s�ϝm�U�c[�A�6! L;����1��+~tC�:�J�����*Pd�? �Ԅ�>ָ���1{˯��0� +�O������B+�Tw�����\YN�髁�g����C������,������:aH��!/,.j��y���b�����I/zȌ�'�۱7M�b����%5Eǹ�ǹy��Ff�[$��>'��DҒM�o��(>��o�/��Z+I�\>K�/�O)��+ȱ�$��W{ �e�\nm8ɿ���E���T(���w��,^ ����h�I�Hgam-!Q��3���e���-,?�~g�{ f`� �Ė���o�?��Z��P��~�Ȑ��aS���bHB#F�N�^�Ȱ�L�E�.����M3LA���`��L {t�"�[B��{�(�n� 
��a�"����]H/�p5\��'�mE�L�uS0��h��`�u�BT��Ŵiٲ�r���Th�1�d�c#�pk:#�&H � E\��\�(�N>0f��?� .o�كOlVÝ;}�5"_m�q���B�ؙ�~��T�a����K�z1S�������Y���y��-�l�֋>���?8��gB�n�D+�cɀ��6iИB<J���[�w*�&dX(���z�g��U��'-��>�f2�.���"������.|����0�0k`�N�	h���ð�������MOO��٢aF�6
���ű��6E��1z|�����?M�络ɀ��O[\f�`�:ۆh9�x�Q�`�g��2�!��}N�4�F:
�:��z_ZzW�콼�yh�ye������n�Y��} +x���T �.ŶhhkG�Đt�^� ���t0->�\{�D�x%��6�@-T>���ewP�����'c�?��//I2���pt*�:���3�K2��(�{pၐY��QI$�X�{��^Ө�}^�t����211�+Ӯ�7�ɝJ>x�����J�G~����C���{A$N�жz^���`gT�cW�����χ�'��(_� �*2r���,��� d�M~��_�<W�Zuf�!kG��zR��uz��5�x�&�O�p����u��ʊ�>)2T���+~��7�� �;�1�z�2Y,(��3��4-Ez�2;!��Ͼކ`�|�Y���C�v���og9��y�s�,uaf ��;�͘c�q�\�Ď��ǂ�$��H�M�Ae�Zq�s��z�꾧���p�U��SV:$@U�쪾��[��Z��ӧ�OC��L_7r������d�����|-��?��{ÿ[�KC||p9����Z#�o�\��	w��:�XV�<�O �f:�j���&�<��L�,�
n����6��K�
+�-Bm�8lϜy���nֈ�.I@NC��;F��W_�a�E_�����dN�Wqr�8��Zq��wvb���֓L�A�mVz��C�H�������#~P�ٽS��;�cY�%��v����T*��$�מ���t��O�Io9�0��{[L�����)Pʐ�q}��������T.���M�i�k������	,����48
�$7��F��&}?��g�`�$Ӈ�N(�3���F?{#	m�&�G�Q�/��w�o�~���
��Q��Er;���1�M�$iiY*K`cm-el�d�Z`�dfG&���uG�2d�,���&�P�ĸ�_��N�Y��A\��`�̘�l����x�z5z.WDDĴI����Q�h(!iPjm�_����@l,HQx��6ĩ�g) ��W@I+)nr��Nj=?=&O�����嗕͘��H��13��0N�B��Us�K0pE�����oya *� ��#�E��N�g������M��e��{&0�H 2���i�N���S�U�fl��^��;aA����ѽZ�DzY�H&��[��h�Íd
�'� .
�R���ihh�P���p|ײ��vj���=Tl �����^�_�͖
�l��wA�>PQg�2l)�rɟv�u8���O+�އ5s�h�:�D\�2,�VE�ۭ���0�V�PN�ل����X��8�&g���iK������uu%7C����XE;Jr��?{�f}յr]=&�z�
�� /0�����W}�L6��� ��q�6~	�А�[|�P�����Jtm���Y��Z|����`�:��.WU�y����V���0�Z%��Ԩ#�\�C#7�������� �v�rc�`�{>56�ӽ��O҆5_�������塚~�|)�����vL?�^��(ϟ��>�Z�I��ٳ�IU|��I,9��%B ֊ҍ�j�ćJ���o�oNM��p"4޾5ӣ9Y�Vaē��gχ9���b��OL��k[�]�uL���n-!L��'S���HK��5�=��=�# q:yT�h4rA������r'��΍��U��l���"�8���!�����9��qN�8�kh?�+���g��K�nԔ,�O���HO_m�~D�����͛-�N��_PP�?^����d3v��y{(���}q̒���ɠ�����c&��z�4$<4�����|L�󔶷��1����2c�[��E����������t��?�қ�n޴,6�G�V-�	�P�0��q�;kI�;����~�f�`���$�Q��\��߹d^��k��K�Q�pU�kkk�\:� ��A��&	1��x�`���&���O����W�Ũq�mMf�֟b�1�(��k��z0�B|���#p�6.�_�=:�i񺠔��G�������A�6⹸����X��6>K��Z�U�K��0�֊�Qgz�&6J�lU���S�L�v\,����dIX�}��=�`������t.�YǙ�� �m
��v�F^[��<�X��Ko�]8�P�Ї�1�1T2M��o|O��1�o�=�BP'j]+��y�`7�T(��T��7qtTT`���rB��^�e�[����P:Z��ckN�_$���.7v�?�^�K��� # �*�:�㕝*����n��N)�܊���֙��I@�6/��^D�:�u��4j%g``�lz�m���!|. ���;���2PV�^�^�C
���!���>�LZOa�A�;p {����ūsJ��� �#>\�Z���PEN���u�<��×�^=�5�g�	*_�M{��^�P��C �0�?�>�Gkyɹ�fM/.Ƭ���'B����2���8����c��3�wGxd��4c>���N)��߼��� ".&����,̩��F��J��<L�"s|��f���l��N���r�_�{{{{��:5[A6p23ix�e���eq�p��w���+�,�Ep'\������A{Δ���:tt�Q�H�� �:~%�Ҏ�!��@�Ѻ��	�?'��_b��IT�N��~J�l��y.����r�B� V�2����" >�ޗ W�t*+�W����z��xC3���R��k�ߚ��A��zl(�R�l��&?�:�!�=Ի�J�'|@ť���nە�'(o)���O�K'"^[�o+'��X�65�}-~�(��@��u��/�텽��L)�O�=��8Oy�ǉ�O���I5ޖ�osLĞ���ݔ���]	@�x!N��b������Yv���"=%��f��E��jI;O@��K#���8�e�;x�p�K��ï
���+q:Yt8�@P�Г!\C��k�R� ���K����p������UW�����ٙ���f�I�uG�11(�(l�0�zyy9C����]�ϟ?zN�@S?�����>ۊ~>	����RB-O���29�����xo���akz�������F��Pk�_ �4��3�f	�qǬG�J����h��1HI�0E�4�X�L.�f�p2�G��&%'�JQ���y���=�U�jط����x]Cø���əX[��	�Ҙ��qt+!A�y��)�Dɪ�1���s�;�_~��N|EJ|^
P����j3i������Y|pLp)�g@|��~
�-�<��>*���)96�Pu8Y8�u�l��A4�׺Uh�Ʋ�g
��D�r���Դ hǭ.UqO�N�?L�;��RC������)��j�Ԑ�Ⱦ���>
"9���d�<�h<�ܱ�p7�*B�jI&�Io@�;�%�:\��$)"a�'&~�fec�6��I��y >��[���p��������H�����?�������F+�;K�	1��M?����c�: �*��?s�s $))M�0_oG�y���ǏZlcTʪ�5�(�5�Z��!�~�#eg`>bW�>Cx���/ڧ��8+˽=��g>T@tgt�h�~+(@�uT����gn�t
	�r~~b��>�u�޽�k���g!���(��^>�Y(��8��t&�<��2�D3B��jI"��W�o�u�����m�f�"��
|<::Zv϶x���j_]�I7M1%�#���ę���DY���ޢ�Y�=R�������������}�+�V=�{%I��=��������J��ᣝ��8���	���t�_�hղh�BX�fpW�[���Gm�I�3ƒ�mr��Y�U��XW����W�� ����N)׬o}��f���X�~����H�K����B�h��0$��R�W��Ot�G[�b��g���؏t�9غ��PX#2���ٗ��\�&�k�J???W�Q�4�����I%�}z���ǒ����v!�Td&���(�F!Z����..|����֑���O���X(I�/i������+�SJ��r�]�?U�wr"a'6�WN��&�H���~��	���\{"���?�����_�:�Y���Җ.����h��a{�ژ��� �y�����옓���mo�䫫)� B��խ�T�όe�>�c�a��vd������ �q��נ!��엫���8�p9DҶ�=f]�6�['8��3D�*��^��=p�/�0�to�㋥|�b%��H���pQGe)P�~���= U�dC ���<񰱱!�[���0ѵ��1��7������-��;2֠�a�ЋɆ�� >��~�A��[���T��jHv��(�c�)�&��KA)�����k$~(�����>lm��6�[����p2Ӂ?������HM.�߿���Cp>�R?�� 7�[��P˚�#��>�]�X���	Ϸ�#��/x����.ӊz�����B�߽:WA�q�aPǮ�q�bwsy<ୂvZq0F~f���'5�����c�B�����I4��?�3'JG̺�[Q�A��a	��)伥n6}ju�V��"��$�kě8S�v�0�vkk�d��?V<���M [NB�Ԋ����͉��;6�v����ǍC����71"�So�ѻw�6^��:��3�I���-�@��K��H����txq�N�sՓ3�p?������r��\/o�
`@icgg7��O���V0F���@� �P4[^_?�t�77���� �4)�����Ծ�ǽ@G{���SS��'�v^��G���.t����B�[�^�@_��|��Y����`���/F�O�Cx3�欢UG�ĥe͞��̴��WaLƢapXX�X$��Q�XNت����)&��eE�é����9���M=T���΍��Iy��`��	A���k��f�i�op�&�Jo��	��F�(qܞ�l��D�8���j�C]:Y)���f8_��L�1;+�/�0vw#�d�����Q�B��ߒ�j�t�$�����tZ�n����{{�/���ǀv"""؍i���7��͑Hp�?.��PJB�j9.`�h;��0%�7* 1GJ�J��Xsb��NƉ�����_wL���1��c�|'_&BU_���,�X֤�FMk�/"/��kt�teD񊚷\��_r�\3� )_��Y�[P0\��5�����rOc�M@�2�� �+���ߖ7G����-�_b����m6�͇��,u�(�ǂV/�����UK��
xA�ݾ3�S��7/	�̬��3zB�,��7���17� ��%��h�iu����ܼ.�:�q�{mB�~/1�@
T���HZ;�E��lt*�<����ĹOJeҴ�\�
�h�!+����=E�����Y���Y��q�sų�&����}�g	ކ܎"vz���3����jfD���5�"ʺ/B����%����d�n:���NL���:
���7����+-���-*hNB�Cpm���
^ 2F~�~����Z�������M$���q�@_'K�H�(��0b�'�Ѿ��|�΢f~rf���z��K��4[�I{���ݓ�co���\�i��!�7mkT[0��@.Ƣ�3eY�N���h)���2�n�,�ǝV�w]�b���0�	�4��`�	Q�����efv6���@l�x��C�U�Eյۡ;�Q���NAZ:E@�a@@JJ:�i)�n�����S������w/?��̙a~{=ϳ����g�U4/�t��e����6X����Ѫ"_�E�KJ�Iu�t�oP�i,�K�Ͳ��#�بʨю��^���t35d��|%~F��[��Ǖ�e���Ҏ?�B\hx3�MdoO<�!ea��)otv�u��ʧ�#;M�l;�,�K����˦�r9%���p+E6� ��1	\9+�Ayt55���o߾���_;�����T�S�9,�4��]fB.���@��Lkn���Xy ��}$�gy"�L�4�pO�of����˹�y!���Bo1��'�����JJ|��!T����#����"�o�*U��l���$�e�G���Y���,�qRĐhB���W��9{�9�@����Ê���.YG�╈],5��;;;��bәb)���?~�E��>4���,����2�ߧ��>�ub��B� ��
cXD�%�E�9�%�3��3L~<c,�	�ktʖ�(��拯��&Ya�A�vO����BV.��H7j+��[�Aʼ��O�[�,��U��ͳXmW����sk���k<����'ξ:��3O`@�`�B֛	��M<����̵H.$�"�^�*���B����rXTʹ�V-���`2&<{�/���l)#�)C��k*�_{َ�g��P �mh�N�&t�S�>��mP��@�����D`hd�82&cd4�s�}���Wx�7�䐐ɦ���i�O<�BN�����
����}i�3]��O��w�NP�W��K[�E` �'�m�M�ˍ�0�}Q{�$(	����S��)O ��Y͸A����$6˧�t�z������@�yv:�$�k�f�&�&I�j���:/����������dz7{J�����������~�i���Eq�E�\�pQ�6�ĺ ���p}��ל���û����V-d��IBA�h��Y��wc�}��؃�V����$OV5�-�2�%m$hW��C�zTQ��1�/�Pl㮛A��G����m�o�	^��^�x]���&�;"�P����X5�8�wO�!� �;CCC��rk�k��TL��r��9���].�-:�j����Z/7��R$)�@���g��U��̳|n�g1��פ����s�,�|r"��wx���*�O-�*��:�c�=[gOΐ�xUPYISm�����>���/tG��U��y�,~�0W�G|�/��*�2D&7>L�c:��lw��iQԲ&+`�\K��]y�ryE��7鯬�YW��WEAc(!ad�(�y�)f��+��`��e�Y�E��P���w���Qըh��E?Ǥ�šwR�8�>��j�E��C����X���Ag�&9�Uߟ+jC�I��z���mQ�V�I}5b��9��v{�����m�����(�go�6n���G�ńk���6���r�Ƴ|��UO��bs�Ȝw�?�/��G)4��
�b,K���o�4q	������J;5Ʀ*�����@��nft$C$i�4|w���29>Nf������5G�a����v����˩�����S5�l>��a%Vr�7��W��dr��[l6��փ5k��J$Ux˚V����߻��H���k�mʂ:8�1x��V@�N��%9�?4C~7K>��f�GV��E�PG���A5$��U~HD�����rE�FUh̛mf!Qy!"�x��IϘ���Cj�Kxr�io�!IY�ɐ��F��D�G����7��<��|m̊3�&�Ѵ1j�b|&*2фpey9���5��K^��E���h�(d��9���р���º�T����c�<�o��$�(Vy�ǘ�++y�nM�^�k��pKR*�[>Y�����Qؙ��>Bx��3�M^�J�=�+��݌�둌�z�����E��R!q��Ҍ[H��i�y����z/� �B)Nc^ � 2@�a��1��=A�(��٬,n�}<�{�����j²d&&&նUm���$����W�3�:J��c!�V��,�6�EI6㻟��X�|�J�a��::� E������6 �:2j���QF�Z����~O�?�5�3�p�mC���]�T�ݔ��Ί���gqJ�����a�އ���_��������C����k��n���P���_�KE�Ҷ6	�G�Fq��3��U&�]h���X7�5�_�ݲ�)���[9��� I�L��d��
p^Y�����!eb�I���"_Q�����,�΁#��w� Lyk�n[Lݬ[y�7F�|�|3�[��P@qL��/������&=[��_?��l`��I2E��'ě*�e�@g��;��m��m���2�K���J����!Q �����kFYN2_n�(Od}��5V�����%�Tп*��^dUc��ȭ���?LR��;�'t�����>U����NV1s�b^�9��v���������Gd0�����j��"ҙ��#z�ȇc]u��s꧗X(1�$$Zlv^�zT��:Hf����~�n�q�Ph����?Un��E�IT��m~�SG�����R����W�n��wC�K��R�q����q֓�� ���Ӕ�k*�b����������A�����qׯ������U���V���v���-)���C�v��m��>��tG2��"F�{��Rbg��:��gL�[���r ](����[�uo������Sb��/�8��r2mlKqÀ�1YT/��^�pzydTT���Wiuӳrx��P��2���>�x�nM1w�b[^Q1z�G���U�~$!'�����9�ALY_{������[�*�fKT��q���M�o�&��n��bw��{�nڲPI�|�n1��3�[�u�.���o�_ܴ2?f�d~*���[t� �D��>M/1@���B	���A>��`���*���}�A!�1��x�|5dgs�Dp@�,��������,��;�}a*'{gg3F(n���9Q�z�B�Q;|��艐�Z�e��-Y��*�T�A+P����m��Q������5����߿⦶ō.c�qc� Ѫ����}#�<*�>[���0lu�4�����٪_��./�����)Oi�ٯ���6[ﱗ�i���hDm�	m*��K�%�,�d��3�,�=��o��m�}�L�D �T�;�*�1�oa��U�����^�hZ)�� ��9�@�����-s��o��2_#q��y�1�����$�4y����{�b��0��Z�7n�x��4���<kr�v���xG�b7���"�B�/�L@>+���#���GN<�D�*Z�)�W�h��?j�8�c�233)�N��F�$�	xZ�AM3}PaH����>�b�����&I��s^);�����.輄�=�U0��y�,�ɪ� o�立��a)�Ksˌג#+uDŗC����� 6�?DZ�m�29%%��^�}�7��^�^e���t�۪YNQʒzz,����U�d�vYC.��RA6����b���  l]�	`��APdh��]�K k'����������i�y����@�sTw��%s���Y�*Ǯ�����I���f����]'@��j���߱u�M���*<��X� �!á�J���Z��HL��Ynt�(�#v
������H�f�LNM]��;�^\��{J�X����w
���}���{���cғ>wt ��Ϗ���=-����1,Z������������7�j_Mܐ?��/<��SZ��,����I��=
����7Ui�@�X��`�U9'_ �{�=yYyH�CU�8$A��76��N��4�9A}�Q�"�q���s 9̙�;�%�OwP��xz���o��]�N���Wa���A<�q����-")s�����v��g��KxO�@�V��f�B�.���Q�s#��:9���.����\�S�Aƨr����g%�������4ȵ%"����7���"3�?j����-�M���wY���y�?�IA�ʕ���苾ڇ��wkg��{+�{��I���~xs�^���~�)�e�;U;;8��:;:�V[�>z��t�<�����+������,�Xm�)GTא�����ӌ׋�qQ|��`fy!�<KA�{���@ӱ�4��"`�7\T�.$�z�T��o��|��SQ1�2�f�N����iR�_�ψ�-��͋>���H�����~0vU�QHD����-,�h� �&�<�+r�V��c.���Px�O)?}�i��*d �qk��-�p�a�V	("s�{J��'�x���kB<�:��@�5t���5��f�����<�?M��\�D!�v|��� ��a�sވ�\�/�ݑ���S4"q�P	)�j�S�N4r��0�����>bu1����~	���GA?� �sD�W}��<~���TA��z��x~�aE������� ��W���mm�$*���/��S��ކ��
 �錏��`4<�&pf�[[;�����ގ9'~�z����pm0n���W�LQ������"�61�W)/k��Բ��:��9`1,��t�D{�U*MRP�C!�k2ﲛ+��N̩q~rV���q��%�(Ѵ�d��=wtw�jrA�c�Ru��) *u�pwFS_�9avt�>��dn�?k%�������]���y�XM_m��Տ&����ϳ�WL�e:3�Y��S�ٖ���A�,t���[D��s���Kq�"���Sn�5rG��9w�ƒ��-%����K(9.Q#�O�.��D罭W��6ӕ؃L���hUV��o�n�X��$3B[�]*��=�Bܪ+mYZ�_�6�b<c�ŁRAQѪ���9��M�"����@w�v�Y&p24Z��M����!���;�bG�Ż
N��W��o��e�b�������3�MM��
3O�G�%i�K������.����z}f�r�U��0Ta_ ��U��ؓf-�Gl�c�'����l\��68���?���%v3V�l(%a�ڂyc{\NE�Ԓ��^�lp�	�Yw��f�Y���ً�l�e ����Wr60�F�i��I��M������Io�K��v`������M�`v���̇���>����_��f$;�p�T�P�1�\���jlg0q�6k��X���&�9���$X��G���Q�KEl~+0�]6�)b���j 7����hKJK���?j��z��RY�*��az�8cpgzH��޶�����Ȅ�آ���Q��*̎���I����AL	{���+>�z�}���r|���ޯ�	#7a����WĿi� ��DuD�!`�j}�B�RQ�?.U�d�@����LlΓi>��⚡�Ƃ�������y7��'�*�F� ���o��%q��? Y�o�����&5N�^]YY�z���+�:$#���,�ϸ��h����د�zߩ�M�2
�v?��+��i˼���F=	
�_}2�g�y�d�������i{�g���\���D�����;�Vػ��k�%e���on4��\)���m����Z������h��6��P)k=M� ��������Dc~QQl��"tK�̯�x���rE��>NW&oФ��2�A�Z&s"�VG�w0� ��� 8pR�AwP՞(&�ӿ��_ۤ@ÁmY��N��2::����s����5L���\u����2��QS?9��˽·S���v{?��[nv��Xgy��A��=��`d,��}$5t���jc���tt3�c���Te(p��)O+He�X�B̗�]���d0�o���a���B`1p���[&��
��V���a��R��k/UU�Z��ᤌ;�X{��e8{�1��{���DE~4�VMM�$������TyM9j�=n��ݥ�ߢX�}��\��_R�sh�ْ= 3�
���9f	��;(��Zm+q�a�m7r��ˮEp�X^\�7y�Do��5��Kuˇ���^B66�Q'��xo�}�#�͟^Cj�!��=����J?�E�o���]ۀ�#���F�I�&a��\$ع�i%��WC3������RI�5]H�e�`Q����z����kb�K=/}}y6xw�h���WSl½�,�����I��lllA���E�(>����yZ�Q~jj�1�w���,H5��f=tuj�{�v7k��h�&TH�l��'����:<×��?���y�ȯ��;�*��Y-)!
�������ТD�a�n���(0$$)�W[�T�>���=��̹�8/M=�e��8�uK�P"N{ �74~�_E2�^��l�>��!4j��|ĲR��B��z[�&��2ss�*a�K������ � ��Ms>��qok˶�E%���U�#����w�]�%��OγWVo��Rw��$�?s;�U��!���sk�����yVE*�I�����..��?
u��0U��o����2��,�����& ���uR��&ft��ԭ�����:D�	�6"d_f!Ý���ܼ�}ie2<�QgV)=���3�)$m�����G�:���&��R��C�[o|�ī�y#�SPrbp�C�����	O�R�CܺKtJ���3�3��5�����U[�4�Gؖ��(�$.h#.Ƌ̖&v�5���s:�$L�≊�N�?{�D��͹/��qy��E�����ތH'��6Ӕ�%����8�	-T����$|�Dܺ��,�����,��" e����SeU���Ln�uә���O��imjV�Ԟ8���v&{�s��x����%��;�J����L�3�����P�x�~��/C���B�&�};����C�N��US�#~���@���S����ߪ�n>�suR�gV��W��a�9E����i�i� �ҪO_噿Y�x]
�7��g �x�u]a���}�z���egwMZZ׎�"��ԏjT��s�s\�>�++t�FFV��c2��;�Z�^:����8c*�,p��S�6h��PZф�V8+q��u�j��D�i���R1��� ;v�%�c�j�����Ԧ�ȯ�T�+��.��!��[�e��ᮽ�W���An^�:����<�-fv��\�	ڗ?1�{zx8 �<�tF�w�U*V�W���h������w��X�"$��s��vٝ+n���g��jy�ʕD��FY�ZQ՞�!kt���w(6azhh�e%��
NZ�=��|AQcͣs������hF0wɐ�#	�A
�q�"�W��@Lp��*%�J��0))il֗�:��T�GjOOS��YI���y��#t��H��I�49��Oߡ{���5X�8C)��f���GR�L�w0q�E�����h���\4q�������`jj$-�/r�rT&S���u��5��A���a��x��4q�ɠ���hn��G��;�|	���7����aJ�s�����'�ݷ�@�6E�S1s�Xbm��/Y����7::��$��������,j0֜�yxP^^��n"�v@�(��wݣ$1$F�V�u�_痮6Sl��_b-n�����!/^J����0Qd�PY��_��]|�]���b
�W5�A��'I�wy��R��J�s��O7U�pcJ��q>�ӿn�B�f�I6���Q�5���\K���%�Q��Q�]��|��F�F�� ��yQ5�Mc �o��gb�����'��qk�ed�sENUY pxZ�a$���G>Q`��}ծZ�"�Ч� Xߥ��P5���q�'�p\@�k���)N���w��Q:=tx��ʶ�w�W._�Xyx��
�C�^�A�HUg?�s�$��"�Ξi�nb��KQ�]�d��"r�-��]�(9!��?'���4%q~oNĚ? ��j+��^\6Ɓ $�"S�5,b�o�r	d��i�x�H&�0��t���0�b��2Gȅ�C��%�7H��`F��6��|���}�ԟHN���ST����L9G`��G�p3X)����j�h�f��n_-((�-���0�?}�e�"�����_��x���W��ͦ蝍��n���lBi�{��qZ�݊gk���i���%��������.���33~z��6y�b�EH����=i(���c~	���t� ��i�%	�Bf��b�[�|�:���݇��t��&7���XT��[��\���(��B�ce]���J+ ƪ�N����S��2�^4�q/�޳���ظ�z���Y�a;Z��'oY�f���퉉��_���~��N��Dǖ�+��g�Ǚ���P��<R{�&v,����C�%KR�l��K�Y�a��tВei�T�����[�����wR&����!J�l+����
X��Q�*�����s�S�c����#`yy�Oi`L���R�
M����V�h�H��Ev�̢�X��!�����m��s��VkuF��	�=c|�-bu4�>�*4y�&QM��DH�>+R[����^KL"^@�Ҏ�_&���U:��G=���]�
�h"����}�O��,��q���~O��Y?4#�9�2L�f?�E���S}�T�	�é~���-���p�1�]����7�"OY�2�᮳ �dZ-
��U�� )4r�ve��!�Ѱ�?	&*/t���8�e�Z<���<�A굱�fNժ�����c��,�|���N�Y>*�-�G&Ӫ�U�y�E��W$g��0& nq�E<��e�ϐط׃�D^�K�T��k=������Y���@�r�A*�^��� �����EJ��;�Å�͊���e��}�_:!�w%�]�gr��.�l
����~T 
�����ی�H��V������'D�ǒ8�V2��!�Y��F0��bm�9��1d���Ox��3-���t�x�U�W](��>H{��*��,}�"C*S�;���.�{y�aܜ����k/H*�|���r��@�KW�9IZ�HV>�"Ǿ������TA���c�#{ۚ�A)�Y��߾Yg�B���uwU;d��M�c��[�h�*�t;�;�M�`�p���S� Y_�!pJ�@��������=*�z���;�� ����q?��nH6U�Gxnn�2�ά���
K�.,��[�T�h�z\�P̻�7��E��k
����s�H��ي1���Z�&%6~��G����x;���[��r�fw��c�ج!!tu91f��JO9��H_?�Z�-Y��|/��[��F,��1]��F.��	���P���!@���I�����n�����ÿ�b����>_���8Yɱ���u�e�]t�l�����f��9Ӳ�"�����P���p�cr����|��Qq�5r�l��{�ƞ���!��+�`�b��6���a	<ß���mf0��r�<�����Ra�t�H�8N����aF(s� }J%�Ye�����60(ׁf������cУJ\��PH��̋$��T妚����k�A�t|.��Q�h���ꕀ��pl��FO���U�f���3�4�����	0�Ҥ �>�B��$9MOG��ϟ��ҧL	Or�9��le���Y�#����3I>9�՚8�	;�����R��3G�u��Z����s��m��aɑ�	F���T���Z o�W���n��}V� ߹o#�J\�j"mk��6�%G���bG�w��J�EFXb��͛v�[@�cng߰ͲE�k	��[v�>��g�}'>�����n�O;vv�|5Q���a�$��Ɠ���RQc4�j�蒱8V��ҀQ�bj�$����4F��5ɹ���Ꞻ�)���/??#���ӧ8N�m1������~.m+��{'�O��8�a�u���M1�N����BSR�=�}�Z~G��-�nӒǓՌ3�;���tP����:��8i��#��uu�,�5�f�3r�Y �Eb7;������B�!�}��N谏Mx6�p�(-$���z�If�G��|�44D�I�@�82�px��m1$�H�Ơ׊�U��3tJ���A�Q�xbW����S6U��8ΎvZ'���o2�������L썋pth(ڬ�@7rd�Px��X����y�J�{�~���3S�:��Z���F[��O59<�;�5���?g[t��o��$S[�r��3#�9��t�>>>��W��zb��J^Sβ0�f�I�$�6�i�:���o�~�Jb��A��~!mg_ ��a�^%M�QuM��F�l	��9��R�.^�V��q+�^��:1�Y����`�z3&.�Mf��Ɨ�����^^���h��R�kܗ�gR,$������P�iƊZuՂ���`��!�
�.���z� �� ���{k�s���^���iD�k�\n�#�������h����{��
�> h���!�<��U4s����2����A7���9�}>_���
x����%����eޓ�:�v/��^D�a.�VUU���O}�0����_�Z��l��U��󋋘��?V��Fv��T��{?N�Z�`�L�<��FO�46O��·�PaT��io�=>>��T$ ������h��\?/Y;�k{q��F>��1��9=��P�eӟ�\B�cY��l�T�h=�]�L�6��ԇ����/W:�8��҇|z�\`���j����yVm��mN�G��Y�ܳ��# (=gEzK��z��z����M��9zV\�>�D�
3 ���N�%���%ϦS�Ģ�'���B�ES�8�ܬz���uu:0���G��������>��I,�/���ާ�'Q��U �jaa�J?�Eݞe2�O0ߡ	�ڗY��Ɵ�,��c�(��#%�xA���+2ss���`�&�c��P�h�(^��6$������������^)>���_���oJ�P��U�a��ˡu,��VԪ�Ǫ+l��9�V��BM��--�0ahh�r�&�o�g;ɋ;�H�~b��ΐH�~*�7/�]zf���gIp
e}����@�L�|���.�)\|�#W�o1>I ��,T��]\Dұ���0����C���v��/y���vUǴ�l�j�~��L��"ɒg�7�0���ec�;�v�+�2��F+F��G�o�m4�]� ���7�����|8ݠll�hى\%&�%�f{�+E��7��Q�N�����dݷ�z�R���2�-�A�
�T�S�(�ϟ��7u�EmY$��]>_Q�t�%Q_q%+/�⮛lu���ڀ0��%�mpe8�C�����k�E�3U޴�|������m����D��A�Pi����Q�'�������ۤj�\�����<�����
"��$̄n�(�fZ�q��2�6�S��L·�.��5`���BjZ���k �jl���o'|4`$y�� NOV��7%1��!�O��~c3℞a.� �
��)�Sⴽ���M��ܷVa�����;kt̘�p����7~����)�/�k���QK��S|%nh��dEr�����ڝ�@���cI2슸���`�FW���k�ܙ�W�>�5�w�x�9�����!�h�s�=�A��~�1w���&��)2r���~��E�=	�(y����uɐ�%*�ʊ|�XI��,�ǧ��=D˯<|�tA�������;ۼPלge�Y�ֶ��P�_�d�}��G����Rµ����[V(�&{r��U5Eؓ��o�8�.f�=,ə�}f�����	�^������i�U�+���A}"_��ns�
K鷬���N9�dQ���層�����wF�����a����U��15�<�mX��l_#t�6�{ϰg�Q!T�e�N[婶K;b�'##����٩�CT0������KnV�{B޼�L�ѐ:��r �ֿ������ݰ��H%�@���8�d�fZ�
P��+Ziܗt�� ��1Y��LG��� ��whoԕs�-}b��%��TN"W�j?nH�	�]��i�SE��~�H��ϥ�����fO�!9��q��x�0�ŗ�+�������>�U������H�ܡ5����cP
��q���lw������2ӆ�B1t�򦥥�m�������S�H)B�p����/0�}�W��	K�&̆;p����& ��a�����}��x-�����
�6��3�^
B��ė���ո0���� ���F�?���@����_iQ�M9]���T＜Bݭ�V(=�˖���4|j�-t���VS��p8��w�a߃��g�M #z^L=���aq,��l+���dw���;m;T����,������;.����a��ϑt{�fA5]_,��n�a�V=�*=�C� ��k�Z	H��Fԓ�(�~��LB߳��\N���
ߪ�~�]�|~�z������W�=Πߑ��e�]�M�~���S;[�����r����$P~�@��f#�*�s:�r0p���Dţ�3�����ʄ*�^��'[�D��N�=�WX�1_�,�y��v42�b���Ț'�Jv��7��8��/���jEV��qO����xL2.444��u������i�M�������Ɏ$��iXt�_�b�H��D..�k#�"p��&�@�F���ݼ���pM��K�����@���c�O��ԧ;�I&8����d
051��P��(�^�Lg˧_�d���1��2�yR�D2B�^'O]�ŗ�/E���GA\{�]g�>~�Yq�Y���f�|�u%���K?�tO��Ǝ������M��~������]Yht����j�v�o�ib3��!I9Py���5��W3��� J�,�:�S�E�U�,�n\K1�ӭ���=���X� m�:}�Iv�W)�]���#�@�E����ox�&����F33��&''u��K�I�+��t\�e47"Ky�˓+Y���j^EB�S���5ٓ���9@lW](��<������%j����Z���q߳���u��Ũ�ҰS�3ޏA�-����;�!��5�k�q%ǟ%���O&z.M"�.}���'�
$Z �A
��1z.��{�Ά� ��*�,Z�@� ��@G�ߧ��aYD�73�͓�)�����˝�.Yww~��nZۨ'_�[�
�j�62YL��CV�%��
��FG���źo����1�--}
�e���!O����r��E��eG���}4�z��b��zgډ_�ɑ�'��T�2H��{^|||��ٓ#_F�R��]p���/�X���#�x�x@�~卮�&3!�Ͷf!)}O{b�Wm7(✇��SR2;�<P���J|Еb�Tr�/� C�QOՇb�N�w�!�<�?� �h��^�^�ġ�sMmcK����(yh�E~��X��*3����b+̉��	�k?��P����N��P��'�'I={F���0��8��!�%F��3�跀�'�w��tٓى,D[\��[�~�ߐ��O)��*�!�h�b9>��sK��V�������y��`�y���k���8������Q�<%�)Wo[N��k�z�����=�[,�В�,,���'��,�\�m>�kO��]WHP0L�������Ϟ;��R�|����&֜?��BE[�,|��PVT�z-fx������p4d��IJ-~�#BӼ�q�n��M��i@�U�]��9����ؐ�����k������sS��������h��m�cc?��j�#����@z��j_Dސ��I�Ƅ�K��	�%Be�\�7} �,4�"FY�X[ki�ag����Xx��-]ʻ[pr/z����94����Ԛ�s�/��L��&3_����T�5_wc�n K�p�N�n���`!7��m��|������mɝp�s�����ߕĔ� I[�89�$R��
1M��ם�gR	��`�a���9ŭ)�j���|��weɋ8�-v�3_���z3��X��NNj@Bۦ���*��`��k�����
��:!E��?�@��\y��v��-�	X�-�/^O�ۿS+��=w����:*4���^&�h�St*'���ziAO��2Se����B�U!'�^g�W<+�%�.�]1��<̃}Y��#/�m0�@�U
�ȭ��q�C�2�w-0#į�ڟw���H�,�k��*�nn�n��U�n�Yf V�'P���'���AA�ԩ܂4���/p
{��\۳�����m�+ZaGd����b����F�-��"����j�'L!R�/���m��g���;ԟ��mj�O^���\b)���ﯢossCx	'O@�d%�jpߊ�,�7��5)�_{�ް�}BGw���B�(�>����{����{@E������0p���]p0v��m��s�
=���e����H ���<&�g�d0�|��%��|d���e1���ON2+���o���l��g�8ȣvŚu�17�tll|Vjq���TUUA�X��#����D}Y�`�t+K�g2�s߿�t=�2��`�������)����:b�	LT�M7D-�}��@�������AR�u��KNn��4��?�%�+��/�y"�P�Bg\�v(�7C,zЙn�dD?{�]W�R��,�PU@H�N(�cE榮 Ӊǧ��`��9-һ���2Ymk^q1Ve�Y��q�D6����rA%ٌ�Q�Pש�����,��B��5��9���^���L.��G��B���d&_����C��J�xye���S�=?����9���|N(�ǘ4��J_͋���X��j��}����w �N�����d�JFFֆ�\k�������!S�I݈���C8�76��ԣYP��`�K���:���q��#V�w��k??c���)O�LZ�ﯩ���ۗ�j�����*\�����"�e�:���a��M��|a��a��t�����2�J�v�>������Q�錰�$^�'�=@L�UV �6�Q|J
٤�0U����bS����^k��ͷ&>��P�������aIN�L934�o>�®/�:3�ɀ���J��y���+�n�hI���Y�2X�����\=��RoZ�i��"=vʫ>���g�GD3��o=:��T�|ܳ_F�q��ez5��Y�@�O�G�����B=�[���X��1��q���]�,#҅"�р�ג��6�F*���ŭYߦ���	
�@$�Q��lؓ�#�ϟ�||�X�?~KG��,\`�j^�2����>��e�c���f�P(�;�E��(�}M��h��¥o�Յ�jY�Y`*��i�<�����A��A��Xv.R�j`"�9�-`JR2n-�{�^�3L����`�\c��)�<$ ���3���n��.���5
��甙�r���%�S�4�cm:a�ԈT�iX�Ȍ/�}�f�������Ĭd$.kA ��$����o���#�n��ō0_�����3j�E{v,F�o�#���ёT��_h�>>L�6���ϊ��|v�}��<�,���{���(?�M�s}<Wv���l`��0!��v��;S\XJW�7�O�&A�>����RT+<A�
�ks0��1~1ɿO&��NV�@kU����^�a�Vl*���I@@` ���Q }y����L__��jxʾ�!��ɔ�WLտr�P�F�1�f��_1��mmlm~H>�E7�@�����$N���U�R�z����_Ljx]�����n���,�]��ʌ�J����쏙�u�Aj�*}x:"ڪu�!/��f�E@ xdh����:2��d� N��!k)����(��������}ˀ�;�w�����M���iy�c]��u_��	�ps��f���w�X���[����%�v��S��ұuT����2$�@�#0]ȹ)㣄|�&b������_���=�~G��0��+!q����{o��q�sӏ$��^�R�?J������,e�Q�T&�6+���l8��`��8l7�:W�l�ً������QM��s�@�uٺ�@}�x~umF�g}�j]P؇	n8ccbV;�v��՝�y�n_��]�Jd+�_�������KC�<,n�[߷9D��X!�B�����NK�*׀Er�y�a���ק j!q�RW�m��-O� ���ei�[�QeM"��?�U\{�����8{g������F3��@	<~<+�����?��"���ׯ�q���4d>��dRZoMܖ���t�������+_�ȿ��J���i�'v��|��<��	�E��6#`�W������D��P�e?�#�Q�f{
���w6K׏�/S/=�~��~3_�*0bM�&2k���ޞ߃�V/��"����`J�ӡX�(cN2_5&C�.�`�<<N@n*���L�=�
Č�1p�h�E�h^ݼ7Z0t*	?os�Ng��G��<��4�����I�cX�����T���3Ѽ����5@�W�"�l�Գ���ɢfϖ�xq9�ӖŰ��N�l-kO'_ ż�k�[��"U�m4��N�X��u�a������| ��(��׾�8յX�aB�G?0�$/�>�涷�&+���C���dD�T���L��c�{���@H�;]R�@��^qj�=4U:�h5�_�������g�4됅v.J������� ��o��o��#a���.��(�����b���#wgj��O�wV�⤜S��e2K[�]�`�7��a�1sZe��1g�۹&���{�)f�N|�jy����"��G^}���b3����&���C�^��lDa8k��**W�|��ު�@�`�&҉83T�k�e�,B��k=ֆFF������6F�����Ͽ��T�Ԁ���A=Y��6���o��@
��C���Gñ+·pN��8ʔ��<�_0i{w��*��㞾�!u��/�>{)���1�T��u��rrU��DU�t��wr~Θ�f����x&�{g��C�O�b�
2@?�J�0N�A�X�^��s��O�]����S��.g����*��������h��B�Y�vv�O_T��;�i������B����0R�I[�o�#C3���0�ɚ�l��n^��5�G8����8콜N���?�P��,�}�������ڸq��L�3ȻW�d�x�)�h犄���#�IDC͠�k���r��jkO� �fEt��6HU��x�M�����exl��3Д��R�@�[�a��l�-Fƌ�q��6�kHZ�s�$����l2+jXntW��n�g�da�c���	]���X��5Ԝ�NE9��s�v���6�o�(�f�x� )�O2--q��ޞӲSS����ɗd9w��7#���UK:���*��7���$����/7a�:d�Q#=u���\o�𴇦<(�щ��,OO��<�=%ȯP�;����:.ʠk�niIi�AB������{�ni	A@��K$V��������y���ta���9W̜33͹�W#֞9N[&����*E��@�8�X��Z��7%j�(+������a��ʸd`n	�̓(����nB��`|>��N��u+q{�3UR4�Õ��%�9�J�x����%!�^<�:lK�?x���(����!�� f�r��:,����o�mn��f�g���D��_�A#bQD��N7���i�y��������x�:�����b%i dzr2Pq�^c�Zf�?����Y���7|�ݩ�/����
�mk�S�þ��}!Q�*of�e�?�P@��~C�E�tۡu��E6�;	�k!j���8�ߧ���Q�g[|��!(�ZA�������s�,�w6��& ������Q����iBޗ?���~<˼��Aq� EV}0�
.�[��<���y$y��Ǿ:�#0(���� ����x�L �l~,4���?�B�bp�N���8@1���-u���5C��/0z^$O�T^�nL�o����n���E(E�����!��	���S/����}l��H���ն�☒�Η�R�N�a�WK�܁���?7�}������#����d&S�)?�,^;�0��#iC��}Y��uI/�efrF���N�NK�R7Y�l����Y^w��@����CQDm� K�6=(>[[�V��y�nӒ�h+�_�8��Ugh$�;��r � ����]9���n�����'[�_��|��U�9z1�V.�$r8p1@z��{���f�E�R��+����;�����\��lV���FxQvpH���P�V(�X��B*cGk!JW:NOU�
-�����n��?���l��Zv�R�E��%:N� �G�>�[�N������O222��b�q����
�X��ܪ�R�?��Y�
�O�ex�Q���^�3Í��\��텼��oSi�ؘ3+��)#f|�\���ڇ��,3����ղ�QbT#��@������N����AV\ύ�����Qdvf`�7�33�`7w�f�~��`���"ٳ#zE�o#�Edp��n����i师.՛�,��yu���0w��/1EhH�'�MU{B�(�<#>=w��N=����^}w	Xj��)�m�!�f�7g��~�u3�U���gY"}���U !�Tmo�>�^�{�G"ܔ鹲�p���	Q�7��I8�R�G��\��NͿ����\������"��ÿjh�ѕ��rH���vԶN!,v��������A��
��9)���.$��@h3G?AO�����2̗9[)S��c;�{!���B0,D��$���w��-�<p���`��`?�`�Mr� ҴA(G�[G�f��i��Q�vE�N��&ť�ϝSߟ{�JU6�I<� ,�Q{ɢ�,��!"̍lZX�T���ݵ�j$nVD��dLT��10e�뢐ب�pī0��_��ȳ�4���fs��&�قT��dҊ��w �G���8Hf��:�A��7sK{�F �	Ʒ�WF��M\K�Qw)A�[qB&:���v�_ld�/��Ǝ'�x�� ���u����C^ڶ(-�� rW7�r;��S��G;�#�B����DDD]��J5WaL1�cT6Z���(=M祒�e���O�cwW��P��?���q����?/�����-�����V/�fcSȊl�逩����S>�����S0�V�� +���`�q#h��o���/06��خ~�l��4H":�@x�T��K�Ѐ����ג�f� ����f�0M�}	�,nٟ�PЏ��(�����X��o�p7ѧ�P����l8�a�x1�J,���v��	�=X��Ђv��L��)����p�KFFb|�F�$���a�j�;��I�9�!qC�\۸�Qs�	[]���3�u��s�Wy��3�|���2�����s�TO�U5)���,��E��<K� �Aؕ?�&���Bq���.
pP��� ���܌>>��B�M�AE�=]�����5�
�vFʘ'ˌ��oO���¢�<�WH�VOFU��D
�
��j��\�u�Ӻ����yk1vRABj�����m��:i��2�`��j���dz_�ت��ֹ����3���ߦ|��:�r��Zcqq�)�n���?!V��M���{J(}ӭ4e�5��m�Jղ+&�,�0`H���/者<7��Z�}�0)Qۋ=���+Uc�����n>�#�6�_�tD<ś3S��#z��2�p�c��·���ד ��I9g���+���a�J�Ah���D3�7_RJ�lgJރ�S7mo�EUII�_q��
���Օ3#c@�Z��]�/b+/<�4i�X̢XSo��h�k�'�*7�Dȣ2�oZ~g���:���&��1�x��j���b���h��%�g� �5��K~[�K�G?��_KI�۬��UQ�^M�fO����f6S�&�]$��C3a�Y��{榛�}2�Eo�M0��=�a�[R:� ��dT/������l���;_?�"-�jN2��������E*l�CJF&�m-���K�Q�0ѫ�3�æ��#�TUUS��e�,~�9������x��#N���봨D/켅�|웜������&6܈��
�ML�G���>�і����T�>�Fq�z؛*ӂ�΅�K�#c}���TaOT���m��K57��$���̛���t���&��y���܁9䚨��ihW�̢���b��~����!s���I�Pr�uj���<�U��g�V�#�D��w�T��=�Vu�GC =P��pbLY3��h��,S���#lT{J,�X��%�����Ma҄�-ɖ�Ӧ+�+3��|�$՟����M�B�Exi��}4*#���d`�ZUr񦣤bs����馘�� ����K^n�����-ڈ�A �S�.���I2�3(�����loۯ��g}�.���NP׿�Y�"�����84�w�o0�"/�j���$���&���-$ue��67=���0���Wg6���e��|p�5�a�p_>f&�Wh�R,UM�X�f�cM'Erp��F��am�Г��A�XiqsíF���Ja<T��p|�T��fC]�~wU?aͮO��l����z�*���%j��hF�>~����ى,q���+��Ϗ��a�gXCf3�!�/��e~9�Dr��ˊ�D���J���M.�p�V�������α��(���3�1I�3�h�1�K]CC��3�ml��뛚���������*1C�T��s�q=�r��Ih�c� ivf����~�B����gl^�]pj*���Č��ۼ?Z�T�W��1�׽|��5��W]_Wq��������Ō����X �:<��˛*a�ozL��L�_2��fL�+ھ�Vv3f �yByjj�2+�錴:FΚ��t���|�}TXs���kǤۨ��<pf�[[0i#�/�P�8����|��o�\����Km919򨃮����-]���� 0�i<	��!yV���E-�/�H �����`�M��
�1��r��C�:q�mV����2�4QO�tś�v�\o��L���]肂.
�Iw��*�	K��S�ݒ�\jR������4��c�mK��K��>����$tY\z�jl��uX/�-HW��u���z(eнѾ�${�� z4+���II�@O�yt�GCdf�f�����º'�V��.$��w1]p��k��h/!���.C7�m��J�FO��^���G2�	�	�#�x����"�M����%+#�'���r���e�=7Vu�2B�4+�y���|�F-�X�E�"��B��d6E-�y�����u��F[�8 h{��7�~�J���E�P��sr�(��"�X6����bw��= ��F.�`���	/��[9���J����[tt�-������}w��B���li����,�ͥ�E��=��5�>Y�nM�X6��C��\B�D�udL�&�D�)F2_�-+d�����-��	<`Nm�ǲ���%8��2�;vgׯ./�g��xy��-)�d��q�{E�A��}-|b5y[�����CG��pi�rh�T�$96$N�@1�ⷚt8G�w㣢e3mWo2�+�/I0ȣʲ��̳=qmmm�k��+��S����z�	!��i\Ɨ��O�4�)"��&����-&
=�8�����(�5�)�o�X�b.T:��i��(C@��ՙ���u�E�Em�4�m���a��T�:<�܊��4�b���b�JJ:q&�E�F"	b�v�+U���J7o�:�|Ӓf��뭡�̈́���B�mY�[.�ށR[��'�Ч+ ��ɠ�Aɵ�~�\ta��H'7#��l*�Ŗ��
�� ���ύ�O~��Jc��vT.]&����M������o�FO�D�e��ߛ6��=�u�[~��=(	���-ӡ^�vm*Y��\ڟ\�i5�����'S��܆aooo,~�C>@ �}�øV�I:]y�f�1'�RrہֳO�p/d5+T���s��r����c��L��k��|o�I2��A���4wr����f��7?�ё���	�O������̜�֓?��;�M\g��a���ō�WhGL�(��I�Z�9�x��[~�vE2����O	U�B�� '��ٶ�ːP�֘�Y�?7y��r�(�ڻǬZQ"/\���?�h�Uk%�ufdf���A���A�ma��j���Aј�8]��z����~wz�O�M�!�w��o�	���"**(�&��:&��%7wp���l�����440"u�������0C��*.��B���ƥ��D�<lh�I��;U���ҋ�Zo/o��A@�Z	��G/�Y�ɞ����-���]��-7�U4g��b����/�5c��:�D�Q?)۸���oB��c�K�����$����	æ����D} &�x���6��3��v��_lҁu9H���B})����]1��©au��}:C��&�&�e��$ųM�'&'��L�ց��V�b��oqA�f;���0S�t,s������韛���VC�����:@����7�|��|�u�/Q`$�X��R.t��b�w�D�T�V��+E�*[�G/̚ϣ 9����sٙ������6E��`yl�u��S��}��D�_dE2??<���<:0Ak�#�����1_:GA:^��d�������N}s�ˋ'�ty5����0cb��`��Ľ�:N2Z</�zrv��E��㱔�	����Q�v�y��ďV��Ź�c�R�pq�\t��v�eMK"Xa�|�� lެ7��d%��wT#�CrֲG1b�8�`�����-�ջ�1�5Ir3�������f�SՅ�$�7y�	dC��f�Z/���m=n)�L���;���r�>v�����f*�g>��C�R�W*7��H`+��n��b�
��b�E����\w�����i]8���+L�i(4�T,<6�T��8,vrwg��y�)��qP��y��GG�]\�ĩ��o�./��D΅O �������St�y_����7���-$1[��H�-@]e�c�ߏ�^L2?���!7:\�S�h�Cj�mx�3Ĩf���q-��R;�f͙*�:UB�}[��gm��e�4t+�WX^��	��>0˩c��fJ-F��my�l�!M�脬22u<�z��3y0���?111�U݂%����E����/b�s�6�(h�ȼ�҇�r��p-z�+?DJR���`�0��P���Pc-��zjVf;ǹ�}�ޤ����W���i��ߨ��up0�(�[�K���dJ�Ƒ�*���)�]��D��툹���͘f3hD��̆���P�p�Z�x^���Y'!
B���n-Q���4B@��^�NՅה��"_~�������F=�������8�M���Z
񯕕�	�zz}�~��<�l��q1KR�J���z�;�Z b�C��:Uc]c���)B�:�Q[�i@<�����Qsf��꘻��;w�vn4|�M��Lu�<��3�^v�go��B2C<L���`�;���c��Pj'�8�����%��S�-������D�t��6�������֏W@B���s)()}������Z��5�C��7�^d-����'�L��Qe�9E��d�P����N��ݽ��d8a��q=�강͏�:p�ϩ=n��B�x�������-I�4����x)f}0�@�U��oTC��y�r0;���x&2��.�Y����f|��g��S�χ�#�m�ޠ֗�r����iKE>ߓw�������آH��s����c�ڪ������N�a����e6����9�����G�Un-��(1"�p��snS�x;w�2�U8�6�}��޻�f����vo�f�y�Z0ڥ�Ѷe*j���f��Խ3�B_�����{<=\Ac�J�p�"v�Ј`C�Hu��$�+>���fs6�N��.��m>sپO�w�[JI�'������!1qW:�MKh����BU��ƣ���O�^,�'s��_?V"���X��6K��M��G��l�I�!1 >M�����p�pꏹ9�ǋ��9�%"Y���c�_���d�}[۷j�VaL�t��L�.cm�Z�Z��Q������]h����_%��^�����ۤ�QUU�S�� $������q�ۻ;��A@��}%�A1�iA�<rX�oqJ)�]�V*Y�L�ܷ�_ǁ�W��+v�_)1!���F�K*�?5-��"�[,*�K���FG��Q�ՠ��2����E�ϒ������܅W&����ִ���m\������ￆ��5��Z�"���Ͱt^j�_h������a����6��ʣ�O��JK��,G��Xg,08z�G���:RU?d�	n=�L�Z���!S|��ZC��!�ښ�w��
����D��֨��κ�Yڋ��ۓص�Eiq�G��X��pv��I*}ܽM�Z�rh�WFU�f(N�\r��:�c���8ߜ�>�X�g^� ��_����h)r��f��i �i�yt}��l2�ܪ�̹�B����դTѱ�u� ��J	.��� cLA�H7�M��B��嵉�IQ=a�nr��,�H$^D6�.�	��Pf��h�y������z=�:w��S;�w�~,N䱉�^_AQ1}D޷8D�þ�60,S�4��~���R^!E%� _���C�7��o�ܤ�b�Wq�����U^� Y �,�ￖ�9]��
�A�˧�@O ��D�&r��9����p��;���n������X\��8����@��燐N��=��@�zďZ�J�[�A|n�HN\���@��8���I,>O���vJ&Z�X�I��=��7/�(9��'o�gN�׍%�Q�G�_]���uT�~|�'���Ϗ\^^��bv6�勛��w����HiY��J���*��PAK aA	�cJ�����(�� �$���2$�/�`H�緵���L�X~=�	���; ����ē�c�8.+_���9�G�&[ȣ�S�h���m��׋�x)�����.��UN<o`p�LZ96	oD���̜�;��{u����v�.UI�!v9�A�����D�,7x\�Y��2� ���f3[�ǪD�{x����_�����>#����/A\�����.���O �"E/��ˍ���*�W_{�GT���f(�������:cJ<��֪e+$�,�ZD��.�Ӊ�Nz�qq����0����%;c<�O-@�~e�c���=���A�]Ψ9��M�n���{e��p�&7�����>��U����~�j����%z��].=;۬�L�*AԾ�s2S�����~��9�awʉ?G��"??'��ѷ��X�]�-���_A��o3��W�.e)		��W|kC&���m���f��xr>]|Xă��=��2ŬO���+ǰ�L�RT-�e����	��lN�e<q�SSS{���e����
s�����7�L�jtt���.�;d�7U�U���}}$	�G�+��2�K�['r3b9�o�Æ�v=?�AG��]�+_Z�wAإJ@!�>�@�|�y���?S�9���L�s/%]ќH�B�-���"��0�\�t�h�%�'xb�_�j\����~Kl���:Jء�n����b���ڻ�?����~ ���;�d@�O�5�D��Ӊ��b��H��N����?:��Q��(J���0��LU���S� 
��=ٹSd��qJճZe2
xQ O�A]���v�M�)\C��G8$<��Ǻ~V..���Ο�C�LU�nTs3��b��F	�b/�yq0��Zfg���y�m)�EQ�Pޓ�I#��H ��V����\�ƈ�����v\ ���np�����ˮ7O܄���kik�QMOO�R���]�ʲ���w9 M�a����w��������3Rѧ����a�<��@��G���R>v�$1�+���g�^�]�D���S��}��
��(�\��Q�������&i���O8 §N.ܝ�V�zl�]E�Lx?S!-:y�.��P�9���(�G3�=.1ymaȂ2QQ�̄��>���!���rڪ]��W���BΒ?HѶB/*�h�!i��"�Яy��FSW������24���%u�#IC�\������I/vp��T�p��-���}A���soh�'�ӗ���_��59������z#�[�P���1�y�)��^a�=ӯ�v�G�ѐ�:���yP���i�b��{��ə7 ޘ(U ����;��ݢ��$���m���p���OSN��Dm!M8ddc���]�#i��c�[��aW����f*���r܋\{�O���SUK#��&G��9G�	080/�R��0�vpAEy�B�3l������Pu��/���WS�+�ej��]�`Q\�X*֊�	0B侇�s��L��s-����,������ /M~w�>�^��i��ݕ��t9 M�de�]T[XXp P}S��	٠��r���G��O	cd;��&7�г� �7и�(�u�_ʌ�v��ĳ�fnm��n�H��.�<宒��L~��;��������A�'\�W冭n/�7�$ဨ�񃀑 3Y�=�*Afe�>T�+�����bx<�s��ȶ����HICt�r��� �\|�kb3|ťh��m\�����WXI��
�.A�A�K��1��j:�Ԩ^Y<!R�*�C[�S�4ih�6��@��|�܀L��}bUz���!c�W���I[\�V��M�K�j�|�h�oA�>�L�����)靁 �Sc ���#�>����2y�3�;/�;�v&�]��)^ZڅMW���I��<~{2�i��,ysU�1�+� =��v���QG`�ķTu�G6��uf�b�@�M>��Y�2�疵�3��A���J�Gq$��YS�]�j�]��J5h ^��d���\Cp��)Ň�E���.�@	��%|r�l1&�N��Ï�B-�?J�.�m4-ol$â�3R�q��{Ϥv:m�����b�,�mX����\�PA I��K�d��`�%޸�U��6�`������F�쫵��n#Z�#���|tZ�BS�S�T��Z�l�}F���׮�dac�s+��o~��z�5�j�L�A������?�,��rkl0ᾙ�OʢQt�p4���۫&"_pƘ>�atlYE��Fg���Fլ����,|���\h�S���fI��k\W�����/�7��P�N�)��`p�����0ɂ�lB�U\m��������ؘ�+�p�>_��9�)��	�K��)A��(��d��_ul0ZR�K�X����7'I1��Dk�S�zK�?.�V��9;t
}3�<Dk��*��t�J($��X��%'*���m$
�N����.@|w�b^ �omi�����s1T&����y���3�!��I^n�0k\�uX���`:??7m�䒣s�����G�J���E�0T�5�J��nRM�w��8�����������ձ\��i��U���Ao/����JIF5�-B����.��q�zÂ����%ݺ����ِ�t a�ĩL�o��o���� _�½!��2)��������᎒�(�vL)���Gi���r�[�������������������������	���6Ϸ:::�K�l�Th��Ri�Ir����bœ��1�����Qs]�Y�8%���<�߰���qPJ�(%9u^��y��\y��S1�)�'Ա�8��q�}�r��$�L ?= ���T#ן�J�<D9l)	H�i�oArf��t�\�K���
��X'����~gN����f�vT�������͝WZ*��*)O#�3ʻ�7�G��ZDD��Ieǅ�`���6~�<`K������L��N2�hs�I�?������	}�&���1F�u�t�(��B�x��0���J��r��0�,���K�K�.�������|�ikm����ؐ݌/�
��%�6�]��kE�4�Mn5"�Q��;x�(�pVT����"����p��j.�ـ�I\����E��L��F�k��o0WO^>��F�H^��#y��cj�c;:==���Y����\���l�w~�%'?���E�FEú4D�I�w��Z�/.�,9�$�+M��ҁ S<A-�Oq-�1���(
Ó��T�@�	����#/���Dc0��S�����uGlׅx�B�xm`�'��O�-zP����H���^O�A��g�j�,�Ᾱ�y�q��_t6�u?�������/ZX/)�|��]·܌��㝚o0�*x�85[MB��	C��5t}�}�^��E���C��R�����gx��۔�S$�vke��U�pÜiH�/�p��滴	gW\շ�d�t�Jqr�|����C�8�ˢ�{�+��9�Avm��ܼ����R蓉�h��]t���w�G��V������ �#YF�C�}��շ�9?t��m�p�u����)���ȱ�}��?�ތ��Ye1N�����t��r����Ȉ��ac1$�nD�C������n�dp��}@o�ˀ�3bi�l�f�:�O�'�[�Q#l�Y)��3��Z����fU�=��c�v9�M9�c��3G�)��n�� ���GIR]���C���Ӄq&��5,ދi����nh�0f��ix�F�M�lɕ__���>�rI죲�z�Df�%W��Y�퍩�@ <rMK~@>9yh>3&g��̓_�v������G� ��K�,<|;䀒]�{|�k&B ~�
Md0[��_�_O+h0�L̹�� ߅c�+���p���c��Z�}Me�⃛@�O0�3�~��4�C,�׿�䦶���c����]�~!@�3NK�X���J��)�_	y�!)��Ī1��W~���/Ȟ� ����V���j/0w�������*g�]�:��!�'�g�f
D�O��@)~������ҙ\Z�U�Y����Y8&���U7���@+*x�ٵ��
Zp��v=n�������z��\���Qe�^��j�FFF��M�� ���Us6M���ʚ�i�Ӹc|���63��s?t�|}|W�.#�sێ?���)k�..8G���X�G�c�[�{��v|���������F)"B���ji9��*�R�^�i�D��f3��KȮ��MMMʹ�%d`p�`D~@�|(s��+s�tY�!U�SK�,	�JB.M�^�1/\ɲI(V����d��:Æ��ga�pʭ���xm>@"UU9x�
��lTҧ���@ Z����066��v!{sjEW���������/������5սXRr�F)+; ���m���o+�t3��J�b ������H��0|��ȓ�R`b�0j.?{��^RQ1��L9��/�u���!��駵	ؤ�pl{&�[A�ӟd��JM��z����{��f�-�/��6&���5�=l\��>�ᑭ�k׌CLl��ğ�_:�k`@�vA- �������N(XvD6-��?�&v�+����G{Ͻ������,�w��KN���nnnK+�@���zWW�l��v�8��Xh�uh]�*�2�"qܙ�LNI1�727G�k�&u�2���jY��!���)hS���߮,�%��p%��J�:�;��������R�κ�hV�v�1�1�ې{��`��7-�Q�R�a.)���)-m���w��ܔ-��]��>[JTmd"���[&��ʊ��̻��.�bE�k�#��0�#���8�����U�X`9�7U�E������f�I:��~�Yޒ�lb�iT���T�%W��]t=q%��ף]��$e��E�rL��ih����d���}*I��[]]�,b����j__S���7��}��'y�Ғ�䗕Y����O	�G�jz/0h�Kݢ�w�n&�l;M��~���[�8�[�f��ʋ�#�ذ�?�xy%w4�t>��A�*���� a����'|ԲϚ�l�;�-�_�F�s��f�R�P-��-%�7d	�̈́�Bƙ�(i!�;I��="��m��8и6��(�h@s�`EV�"+���)��mg���p%�k��r*}���
�J���;<䆛�i�M� ��~��O"ek�{�4����qQ���
s0�(ÞF0�A---�1�\i��{MY?EC�b��ݾ�?����3痗t�ud�S+��}j���\h0��>�����_6�C�໿�1<u&$$, #�P�����ֶ_�wQ�{t���X~I��qi���, �#��;�I1��}��y*!4n�0Ѯ\����ͯ��&*���PC�goo���頦��S7ڴ,i))�O\��@���Ҳ`�.�$F����띹�����{��dzlC�_��s�&.����Mq�jCb���	�\[�"�9�R���ӵ��&���2W/ߡ5'mr(( ;��K,��y{��g�cm��6;����)L3��~���k{^��E;��J2T�#��Կ`H�$"�^��vGp��ow
V�F��1�j���_���nT)o��3 �'w��C?��].��	p:���+z�������3�#��������"�	�i��v� ݠ���s-�:�sq_�L3T:{C���_m��3TӶ��40����6�� \@d$��{~Gy&���C��{Se��4O%����#�?�`��}��f*f�!:I�Z�}���鸊�摑��<ZT��G@ �6;��2?��i�M��kl\%�X>6d�l���t�8"+ЩjX��/ �V�)�\��q�o�o&{Δ��h��N����_v��<?���׿�i�<�M6�;���;�\NX��_��PٳZ�[��hJ�M�e�¦
7�;�2vh흰#�L�K8tJJ�]M0�{���Od���u���e����dƄquqYI�ȑݿa&@ H�OL[~>�B���o��B�!��8��e����h�J���)�N��K�灶���StT4���:��aj��9!��*�6�{	Aw�32H`D_c���9��:���j\�l:5W����(�N��n��qGGG�����+�B�b{' g��3��a��#�^�B�����@��o>�ЃζF�*�x2�xE����=�#�����x} ơY��,���uV|��	嵔
���6�NA��N�?�gy�������i� ξ0���eA�v�����W�O��/xQV��A���>"�=p:��
	��y�)?�(ι鮭��C����!����3�~�X����֯���רڽD&R3�hMI��>�»�y��v�o�9�V'�ҔeD�|���4�&K���3�l>�nGwG?��ĸHa�� �O�� ��־7B�s"�1�,R�"�G�77��F�B>���4�����fx��� I���&w����`�_k�gj�۽�tFPPw���`��Ǐ��_���|}}��)�����o���>�V��3�Q����.�?U���q�R99�Ţ�M�6�%P�n�+����,--�N��![�N�?�ᶺ�t>��񅆅�` ��ͨ��{��i�{PaЦgsɡȎ����z#�&+e�L�ˤ��F����۱���ܥ���_���8��J͈��+�6�����O�����un���G;���<���0�)��U'ſ�"���n,�xA�h���P$�i����b�SC�]d���V��qP$��9l�;Ƞ�Iæ?��O��p����rr%�������^a�t��BGZ�N��^��L��f:.��e���0��L%lC�J@1�Vj��Nuai�Z^n��܎w�!���Κ�?0Z�u�@�.���.���g!R�3Qǝ�Ke:,��5^:��$��(�Q��F؆O�3����l]G��oyV�[ZH�� nN�`-��\lu/���'�f�I���Z����������N�7}���B��R)��s�t��#��v]b����N,?�����c�:�g0�%0��Gb�u�п�ͭ~��ը�L�S9C|���pv��Q}\�\Pw��]`A�wS48�giJ:M�b'�N_#�׷ۂ�1��L��U���� ���g�u�Lf���Ps�#C���n�BLlƙ��[��P��g�zs&��z�Y�[#�H���B*ŨF��Q�|�c;We�r���DO�Cy��x3H#+������AЎTT\L)�t�5Hԛʢ�0��8��<)�`���Z=:Y\RR0���jR�� ��ړ�U����Z�sK��`�x�!Z��ëI�Sv�uz��rp���J0�X�W���WVQ���� �-̆SPZ�V^^�Ns�1�l` ��O�*A
�M��b�}�ƈ�^�����ӏ�Ŀ&J�䇼
/�E�L%@Ps��4~VBP�pu�����3���Rl��u���]���r��0E?�m�JǑc%4mo�r�}3��^��e�A�[�E�+��W�#̼����J�d~�k��/��������H�X� P=r s0�yUU�ִ)������ɨ	��9wT����]GHII)�&�y=AE�!�ٚ/'�"d�P�[��n���vZ�0�0]�)^e��}�hAA�5tY^����1�wU�����ZX�pq�����|�k;�*ho�����fNV|4�T	��B'��ZS<`�u�Q�x�t�&�+�4ц�x\#��/����^��zкR�d^s3ߪ�����3G���,�Zr"$(d����xe����5���^�݊S3n���Am+&�[sM�19"�}�� �!���e�/�C���Zx�/����М��ta܇1��{������ �CCyH����;lH8-2q��u��
���[m)]b�)���Q����M ���#P2�#Q�wك68��D�ϥ���*	���_C�д���[j �y_WW�5/�x�@dR��b��� �}_y�R�OG8=tt,LL����כ����I���p$���i�a#���P^!���Ғ� ��_�2��`^�А&�-f�ｽ.��+筕�T��-MbM�L���KY[3�2w�H�A�ϕf'ҫ;�� ��M��l�wo ����o}�Z�X�G�tv
z���H��ʀ�O4�h��T�� ҌG%�r*c�ܼ��RRRo��GG�Vj\�z�ׇ`n�6�n�`�k����, h[T�xlqNk��g�����{�4���!wB��y�!�0R~�Fy�}@`(q��G���3A�lNK�����Lhh��g}�đ_�S�11��?WR5�i=??�,WD�:�uO9��;��D��a��:�̹H�O��!��H�b`��H��(�@lu�Ȳ꛷�kk�K���ͻy:�ㆇe�45-�[�9���޼��g��q��r�.����������$����w�W�<�_�*��
ev�0����b�'��� e<�[��w�ᠷu���`@����@����\baV�lmYܠ�R3�%��#ha��ֺ/�������	^�G!��	Y�l����D�;~�_�i��\�#���� ��qeM�q�Ր-�K��ph�>�T���v��p"D�����e���}1�*zm59�@X [��AS(Xm���J���*�.��tl��]�5�n;͗x��y	Ŀ<`l��#�e) G;�2!=8�D�0�8ർ����q�ߎ�p^�R:�T�����d�x���h�kE:pa���L��q��� ~z���D��'*�?��ħ'CJ;s�O����َ�ڈ�J�m5�I\~�k����Y�&�<�q����VT�,
�h���[�Ǝ�!��ss��\o[��u.����2�һ�P2��ޜ%�7!�+ �����GW�KjqM��6A��^o�|)Y`m�i
�a�L����V�M�0 i������X��{�0�K M�LsqEN��l?�9y�����n&wn[�@��
�wKa �������V��O#��\���4�leV;������<�D�����y�F�[6QYS3���q�>
V>l�C�N�����Q��Dr��i��7yqԂoë�;�����z,,,��a����l�g�^%� ����GG��z7�J�����r�/H5��QM0�Zɀ駪�:�!�;�708�D��4^�,�K�J�i>���J����+ʹ�3��3��KM.�������hZ�0��/Y���zvzG���Hچ����ԟHql'>���ڒ���^^^�a�ܳJ�����ӗR*������zuQ'�W|�3�wU&:_�%^����|�vT��.�;m ��a��_��er)g�nnnZ�ۇ-�rv����e��l"���m��^ER��(�$�(���jG���hY�Tn8��B7�w��]z����Λ��t,@����Ay��·i3k�ɟg�Э�f�~ �e�d��,Qy���.�e���n�Ly0@��]��:�Ȫ�:%.Z`��t��&щ3M/(�b���1��;)����E�d�D��e��F�V��{`~�̈��G��f��s���_�*#�q�n�m/����lbܦ�iAT��y~yG\��]R���\���5� �;�ٿ�o��� :�fhiҰWf��K�vvf�ZP�kb8��vH>�]��0��4l��-=�HNM��T�<K��p�3��i7�S��1~�w�[��`�cx�0��"��>C���-��U����QM|���4�WB��~I"gM�;��n\�S�~����
�8�����m��\��C� !H������-x���{��5����������֚E��g���ޟTUW�����-;44PSS3q0�t��:jv�Ò����r�1؆���I�oi3��Ʋ !�Z�2"8��>hll,hg�����p���G�����Z�AQ����Ϸ�T<8��}�P�1=��&(x��r�{�u�MC�>Q���)����XYm}�e��״��`� ����l=�H��m�7{��_bp��C�A��x� �tS�׍b?r��5V���-�Z_(�Z#�}�5��9�$M��h>�+�L�)yN]���l~$�YmT��T��+հ1?@p��
o�g��M�
O���|������s������QdT���~����ݐ�g�=BL�.�~}�C�Ռͫ��0Ǡ̌�͕����rK3�66J� �
��cM\�Q�,G�oH>Ȑ#���#e�D��̬ۨ���@�Ȅ�q=�5P�!�)�p���8�;�6�k�!�oM���r��$54p���S|�ڛ�����f�SH1�:D{ �[�t��Y��u���Q�e����c�����vij+�Cc�wT>�bi�VZ*5}��;�C�RI�!S���_,��𚆧��4�@��UȠ�����*�l E:ͯ�aŃ�u��ʴ`�蠸���m���ƒj�����qg͉���0"�g%�S��?E�ި�2i!��Tٮ
/9��~��S��ښ��8�Dc�_4�w�E�4�A��+ǃ�g�ப�an�;�L�$��d��r����+H/֢m�.'�$��	dn��ݽ������v�����XT �P�A�r��}�֯ϴ
bk��*���*GT� E��ߐ�~5�i?O��������r�0c�tȞ/@<�RR���0O�9}�����|��#J�ғ�+�TP+�z���)M>���T�}���#i����_s$��Z�i �d�uT7�-E &�m?�"�V����(�?<�~�|��mp�%<�^��^x'� c�C�|KY����>&
B��Lq�Kʤ����#�/�����Y�9�4Quuu�22T�G
�߾��5Z\L��@;�m���-��I�+""�$*��B z��Lq`���냺�7����&�2O?�p����L����o%I�:I��Â�"�Gl{�+3��i��CzPQQ�u�E����*Z����&���Ĝ�8����\/G�'�0{�����y͔�D��a�	���T��}������_����a��<����H37 Juk��.gזe�ۻس�+ͪ4!4v�PǸ3������.T5ӟ\会,	���v�V	�rܯlǦ�������h�G�ϳE*5_.���Z����� ��u��hB��3���?� ��k5����*��?d����L�Ĉ��Wu�S̻�>(�/=T�pM���T ��\^��j��{��Nvmj~K��~���~b[]��ݰ�#�����fN\���I�6a%���UQ��k�ֲ �j�o~�{߄����1�ɫ$J	�%vy�J���i2�tu�QT�������o�]7�uv���s�r���gl�������]�����xb�珨���:�ٝO3<~z$^a�Rmil�n�1�Ǚ�u�c�e"-m�G���	�⧻�l��U�5s}�fk�9�� ��~�8�����Si��F577�D�Y�	�߽�0�덭*��t��_�*����S��C5���bRܥ0!���Fi<:���9�����+�1��2��͢dj|��)ͤf���l�f Gd��r�>����L�F��'o~g�=[�c�I���!�zx���п��^[_'����XxHϵ����2���ľo���ZҺ����m߿O��Rݾ�c̺\U�вg�����|jHf� ���ed*�ǺjQ]���'�q*��`��RQ�#d����p���#��# ��ZZ����muF9��P4���YX�MLh�N��u�YYY��_o4�لS&E�^)p0�l����N�ò��8��S�kd��d��}{���쵁���*�u���F���Ʃ�;2�#`B?7w
N���QS	))8@#:R���|i�Q��o�|�)�O�~u�_Ad�x'��`�r�Ntr"lY��L�(7@�b�"Rh})�C���FDn,����ov��w�|p�ܲ�.:��?�"9��a!5��=�������<����U�o���m�M&�zeee*0���,�,��]ʊ�xQ�#���Br�x�_罦f�,uB������R���G���='CCCʽ��l���H;��!�4 ?W{佉;T����>�l�m����Bmm�ݖ
��Q�Jݽn����ۊ{ɮ�o=�� �O�Q��u��6$�v���o���xI~,EҺ�Cv�\^�njj
Z��<�Wڽy�����5?�U�� ��yF�膑V�;��\�Y����7^����~qt����kY�Oՙ���+H���"Z�`H�2�MHL� ��楖X��*��5a���Y�0L@�c��.�YP�x����\�D�֯��|F��|�(�U9�o�f]R�pg-�M�~ �1��!PYl�������}°kj���� ��ų+I�`L�8��C�5��f���c��t����g@(��ңM/���uI�������R��H ����M2Nv��}�ڌƧ��ϣ���ʫ�@����"}������2���ީ
i�´�a|�=�Z� 9���oafX9d��LI,����f;�K�����ǛM���*{q�9 =���xnoh�s����QS���D¢�"zF��R���H�U�iEm\���O��G?f됿;���$�xY��b~O:i�AG���|ú��{���4�x�Ȼ��q��U�0.A��Nm���}}}��=sɟsé� ena� HU�������}�i�يͱ�l��>�9-н��3�B��w��+	�eb(�{XuA\�v�92��3�0�~Jɢof�t���Y�v<����	�Z��sm1�qT����eͥ��l�(.���ێ�����n��*���T;�b�''gѹ��+�f�gƷ��.��}�frb�GYU5�ʌwO�]����z1*<..�+����o޼�������l%Ad ��Ʃ�U��c�F?��@��}�=���W��|�5=a#�����91�����V�J^r[W�����Mdi=A����'" +����f``���� ��j���x.�V���*���>G���A���{l�X��nǔ�qV�c�t�3|i�S�w<�S��-C�ܲm$G�������5׮�!9�6=�$��:��.}Quu���2LTxv!�h 3�&�L��p21IjiB�i�0K�ަ����/�jO8���R�{�� }����-�e�BS����°�$q3v�BEJ����C݌)α�;Y@:�tGRM�`��p����y�s�5(&�%(urZ�qd�/5�" ���h+�Ã8ν�=��B}�L��8��<	�m���B�wz��f��pr�в��@��[��͛���n 9]\��b���C7d?�83/���E���׸�[.�l���������5)�otD�a%���G�)֪�5�PLY������䉺�k���A ^^]���S�}*����g`��ma��	�2*&@oCu���9������X�\\���u���� �Е�K��������'q۟M��[�� �J鈙{`�؞�|�eP�~�!`�{j&$�B>������ 7��*V�|����^�e�1Z	��d@)�B*�
7�z�ܪΙ9
�Y, ����cb�++1"�{�[U��*���P%��Qi�[���7`4��9���<���F���5���똣}K#C�M��v Ͳ&7j���fc༿�l�?]�="��9Ʃw��pjՔ��Rn�,���:+�=o��OmװҹȶM'�Rb��'�)�IZ#ү�6��;�b�蝦;�؁'Qi�Ln���^�n�x�J � )���X�85А�����~{�:�ħvP�*g��>�p�&q�jz�t��Q�r�54���+�3��tY�@)1;mv��ۑ�9���%%�||��})(*~w{%�*ή�}�\l���͏�V||H�����oSY(H��|��M�=��]���z�v���RfP���ņT*�"�qܷ�oqyݶ4:mU��z#������v��~����H(���[Ι����,�[/����;�a��u�*�w�ށ2GC��M�Ӂ�ZY�SPVfm���Yy|�`$;}�����#퐸�p� ��6��/���K��dr�f=���J��8�d0f�v�Fd�:��ߤ�yw�<��Z*���-��<����F���_)�����q�Cߨ��i�g�c �J�p���?I�,E��xc��Ν�"wHRb)�%�DSL�G(��9�h;��B�>����1��$�xxy?~�u�:���T`���ݥo]�i6!�~[�ef���)2$j6�W�����'?�"�����\�6 �q��:�|�Ց?���	�S���J21��ƒm��JpXR-�;|:|�DH��Q	�+��h2�omo��h~��؊��OY�����wL�%q+�E�լ�WM-Ä�o��ڛڡ�G���.��Mϓ��_6Cٞ%nCY}�ȟ'B'��k�s���I���Cy��٘��ʇ�@k�+\�ͳΝ������
LD�R� ��
IQ�M:�{{b���溿z��^HCD�`�]h��ma9�e�E�Zd"��:����Q;$	�?�LW%�PN����'D/�u�ۦ�nf�AY�-u���\#+���b%)!��m�B�k&�!&�o\�b��g!���屍uSȶ�PJ�ׄ�āS{�jj8�P/eT�����<@w	�Zȵ��T�: ��.�z�s)�w/
��h�4HO@m]��%S.�2�s�UUU4�"bF�>{e=at�y�\��Q��~���q4vpy�>��J3!N�������nJ�&���⾾"�.-�c�Q���,e|$�=Wc/�tH��A� �+z��T�W���F�KMG��8s���Jt����2R�<=	��L�#Þ��؆� ��2�f�j�c~��`�{���ze}�j�Bz�v:n��k�}���s�wvv���p����9�WA%Ij.9�y�jl9K�62;*�^z���r�n��pἽ������IQ�X�����x�`#�[?��~�?�2K�s���d����`���ĶY�È���:۞���i/�6|ꋓ����Tj|������×] i �/)@ġ���z�P ƚY]NB���6�H_߽E^Mg����|oHw~� Bh�?1��p!)r���������&<)(#�g�gO�:��M-��^Cv%��m�U�_K�b_�����`A
%�C�X
yx��d1���uﻎ�F�ZY�ߏ��	ԧP�� j�M� �����v��W��A�<CD�ߐ�nl�w�tnsG6[�d�ʹWJ�i�Dx큁�����+�;l��^k4����������
c��d̫uҹ���#�ӑ��_Eo_��4�4H�NMM��ZLXk��/���ļǅ����eϥ��������ݣ#���i���?���~Ki���c���Q�H�㋀O��廪�~\�Ý���^�� <͸ �X�
$xcz*8�%@y�:a}�433#�y, ��p�"���nx�7��Bw��q��so�{�<?=�$�(f�= T��|�ř��������9�&Y�);?wz��?�#����u	�Ə��y�KHo��H��v���V��v�(֯y+8��lhk��~C�f��R��^>��FrQ6u�GM9����8۽������NTT5ZC���A�n�e�8��#Ԑ������!��x�{4
)}�	���R�!s[�Ĭ��0Y,B�rn���;���:��d�v��!cq=��Ǘ(������	j 	Cɕ�u�xvQH�M ��/]���DJ�+���C��e,���� FӘưj>W���n��6l�����G"���Y�T�lr>��4] 8��$�Т�����n�V!2X}s���8<�F3�&�lu�t�u2��@���}Ȇlk7����Ϭ�HCm����0Ʉ��ev2W�*9*ܳPv�Ug*.1�Ŕ.���5y'Hc�FP�gG&�r�=2ĥvg�R6�{�M�V��1Q}��ʢ��B ���͋�ӓ�l֏�]=-��D�"縋�T1��Pl$���C��[�*ZN��6[b��JrsN��>�M��ٵ���{ N�FxTl,k[;y�t�� U���Ⳣ�-ch�Wy'��LP�+_\��ZӤ�c�.%�ܜee��)Ťs�[��9@�f-�^kK$e�6�U?��G��&%`�������D��!��Ʃ�x&ͪq�D�W8��0c�v��f�r�r�Ѥ��~��v��T	;��&t�������Z�Z�e9�f+�49�u��H4���eZ�6j�5�.������Gpt��
oἏ��zB�[�W#roܞ�&��|NNN>�t�:�����J+�Å���۹�e�멹������)7ph��0�-gʴx�g�F���Z��"Q'B�8S�&�|mNC�v��#lrrR��6B�������N���`Շ+����6�L[��i�D�S:ߩR�_�#�4�j2�^���y���{B�@��'��/�kMz q�1t��	�u��竌f ���/���)5_nÊ#ɡ�_6��I����#"����ɸ���J�lƸ�浇��nI�X������{�%Y����K�d�����g�x�&f����.�v(~�e��4%���,�@vT����x��}]@^\����{r"�*N��aww.c":��|6po��}εu��� ([o�u"'��X}r8K�1��<u����~�:�]�|yd��M��g426��1��L�(�\��é���{����Q֝�Q�S��o����s�ٞYc1���@;5 _)S��WGZ �����W7�ϻNo��9��d�=��l]X�R 9�A�@�+�t*�R6#�s�sh:�%
�v#_��@=�ʓ�<^2HR�=HQbAV!�<�>2�S�s�o+��\���냀tC���1�fl.T�풄�hv`,�Ւ5� ]���?��7K�V�~��κxܷ����8�I�K���	LD�]�h]Q��=�-��=��˽���c�s/��KB��C���g���?4
J��c��"�o9vƂX�%�>�ޜ�'�=>������DKC~��A�a�0H4A����l���l���#=Qc1TGn��%���~cV�U^0�i����o��x&ͼ�{� ғ����t�Jғe;9U2����'��,x���	�`J8�xqmAR���NPKr��ײ���h}�Pbp��\�������*dGe9׫�'.����		}7�_0jXĊ��J��g[_7 ҹ��n5^.�͇u�9|A��X}�h�3�+f|]d�D4�ߙ���'��z��om;1���oH���X+��"����;U A+�u�%�����. �$w��-3�5�'(��=H3���^�R*�����
���f�:k�G���/j��d}ʾ�SA���y�����i ݠ�������#� \^]1{f'��Fw@�*N�w�~�KkZ�]w��p���@���C��C�a&>(_�����>7:�d���ȵ�@��^cK����K���,���;	��Y�W��$x�����9�����3o�F�Ԟ0U3�x
���9��&��k���F�2r��}(x��vJ�I@҂|_7�$�Y8��P�N��;�n�C@�n��L�\��m:�@݃�����&��ӓBH�Jr�7�$��l\\A���n�947�Dȧ��܂ܪ�����
FQ]�fEׯ�C�������IE߅i\�o<��*Q� 8��D��R�Ѷ1X�.�>��s��PbtK�[<�FU����@���.ϋO:��F�R�l�� �|�c��9H
�6��r3I�Q��*x� {����.v�jj��"c �����3�q�B����2h���s�n�#��P�!ЃU�FA��[=����[J\2�|+$�J��9{2*L:���B��O���B��KjC;�zρW���	ߓHזp`�>�!�Ѯ2���X泻W����u����R/�����7IO�ȯ��'ޖw��d��}{���G��8�6@��!TĢ��H$�~��S���sBb���l%�BJ�8rWjK��:�Q��pZE�� ��'��Ԏ���m���o��Q�r���ң(Hq@ۧ���%���C���$À���X]�0F0��D9�y�:p*��1��@�F���hq\`�!P1O��*�椠���Sj?��קp��xR]�/��i
�Bk�1�%����rTPV�����ϟ?)K/�Mn���:�>i��4t�!�wQj��O@���1~k��;��Q���y/�����&;3���gLx�!�P=!@�Q�QY.���ZX>�6��:o�N��AƖguH��M�ߠ��p��CyB�@~����Y�_�&�zr��۸'�;�}q舦��zt
�:�@�&1@�?����w���^�H?�!X�Q�p�'�-�+������p&\ �@|�ME�\Ջ0r��Eh���s5D�l����:VV�����Vip/��t��v7�r��y���	Z��74X�/'}��YW%�@r�
��0+��w_l�Z��O]��7a,��bH�$'p㓬��|�j"ݣ�$�7�̋�:�s���xxx &ym.��$$�rP�Gvm;t�9s�'��U�+�{5yNE��� �Tj��c���Pל�*\�1���� ��]>�<�k�t�yxV��k���_��`�����'�ߗvoۏ�|�@��-B��A(@��y����ls��l)�z׼F�[���&�I'����%S����?�A����fB�cBp�4�zF.0�Ho�]��/;:2GM�� ���2�&&���5�9�ʴ�V]�
a�����O}�R<]x���J/��ȴ���G{4J.���<!��;�{gvr�Y�ͱ��W����A'xs_�����Q��/���p#Ĩb%l��m:V��R���u�e���!<�?�&7��~T!S�Svٟ�z��R|P'����A�>�}��ˏؤ'#J��ʔ�K���]WnE8-����.h阾���2W�E-mF�V��Dè��d�rm[��x3#6�#H�X�P����0U{
S���%�f���)�z\J|�@�F��B�2����1z|\h��9N�R*k.- �!�#��a$2����s Y!�G{��2���t�rs�Wεx!x�uO����l�F�<Y�+Qb�m������N(D��춺+�a�y̲�����9j�f/)M�L���-%#)
��A�,)#��O�G�=e|�]ZQV#xB>�ǟP�Z�1���[��������:s#(3�^:� �����h�Ԏ�;�۲U��-�nD���UZ;_s��ŧ0帻�c���=_w�o���<�����sʘ����Oϙ9�Y�؉����K1ضs�>:%��X������d���5��٧�8]������@��8/���K�r<�����WN��y�����>���q����/u�M�JX����#bG���0"�ow�0#	X���c6����Z���,5���n��O�iF�y�@,��iӉ�V�!���w��$c�k��L�3K��c��t�ي�F66����k���|���}G �T��Q��"�7D"+�"�,6 R����U}?��q�����[��oé�l/�hWY@a�p�݇@�<\w�Y�"ԗ��*6���3���7
�;e�ڮb�m��0�7a�o;5NZ/�^�^���h�/À��(��<�8�~���4\��B�Bz\W�н�n9i_�(T�k:��hk״O:E����t=�~�	����	FZ����iNEh'�V;m�_��j�w�
�P^^�z���|���@�:��v�U��v�]ߥ�+Ъ%��b��	{�����9��<����nM<�}~�=�D�%%����e�0�%V�����Nkr[�G|�Y/۞w�B���7�����&�����(�T��8|OR�9��~UmM,C�U^����ol��mn��
V�n�d���*<�
�%J�h�)}��'f��{�� l���D�a��;�#��%7�~�ngj���vv����`������ͼ6%���*���s,$�v���-���ڸ��`|�=Я���o��]�l+�������>7%~�f�a��R�q)nl�����q-}�ef�����m^Œ_�4HP��	���^v]}b���/�[�-JB�"�{r��r]��c���Gf`<Ht뺅B۬\�C7s�B�AF��U����*Ha�cq���ܚ��'���ˍY������/	��U�vO`����x]s�[ܕ�D��r/��KK�9323�ݵ��H���^ƚtЁ� �K�[�9�G-�az�F(��2�/R8au,��g��>��u��n0��5^��	��h��ֳ�GM:��.G��g�й��,�E�~�����U��lSn	UKE$��I\P�g�e���+�s}x1��U��iで+�L�5g4T�n�G}R�ͤ��Ud*�r�~�߁2�����U.��XZ	�z>���Ru� yG�Ą/��#����ؽ�^tad����gi��[��ۍ�(vߕTOl
ؑb8�����ǣ��O�-�ڕ�_9�OGC\�_tB^�o^��_![g�>cvЊvq�7z�gM��J\��Z�AN�=������-.YK�ZV1�G���;w4<��?�9��i��#�bo��	�°g>i��_�-��w2y����t4�@#�'m����H��s�>�E,Y�S�L��K�J��*�c ��D>3T_��***�
��W8�c`2)޳"�@���n��-�Md�������Y1&��̌������g�͖B��;���n��:M�o&�>�sp(�~��@
�����_�z.y�{ Y�X�	�䠲�њ����FY���FՒ;A��#2�J���Mda����5�w7��5�$000�GGR���:��nή�F�?��Qf@�Q;���OU�����{bƱ'�Y��]�|�V���Ό���,��j4	C��?2��*%"$�;s*�a�)�ؗ�G�>��	��e�C\��R�s�=�RI(P�]N�z˽m��_5����D����:�>/�uf?��{BQ�����E-a<�6��>��?�?��u|�9Z����=a_}���}% ��^��>#�f@���%�1�3�rv���QXQ�,$��fe@^�W1{�>5Hcٹ�BT���P!;p�3 �i\�V��"=��P:�3IT#D\\\_**Ї��)Y��D|k_l~[���


Ԑ�����"H]b���e>gp�"P�d3��mF]S�z���Y�U��gE.kNA��+�v����ZV&Α.I�v�(e���BDDMR<e�� �p```�pi��
��o-�o��Ym-/�V" ��:�����X�'�O�J�F����Eb&+����/A&�����**��31)L��CH��w2x�ɩ����v�#��؎ε!�җ%v$�HI,k]h��Ob��� �s��E��S��=R���ԯ7�R����������\�x7�cE_�^E�߾��������y�F��o���
��I0	��6j *�Ϭ��ef#���ׇM[����p�SL�C�2�u�m��>z���#r��c���T�y��29�nb��+H���A��in柞���G�#�*L�`p�LJ�7?���e���UӉ�1Ϟ��R����]c�BY���,	�f㼺`�dm��Ey\ұ����]�gXpQ��E0fX�!�������Mk�8�ƒ|��L8Q�� v�xд�_�?��fQ�3�m���<���LJ�;�|�1��o �~��5���8/v�z���x\������S��O���L翿��������
b*:;A�xd��Ĵ��nU&����!��w����_���4k�M{&��#}��Cs��x'�p��m�Lyfc�=Yȥ�r��.����[��?Gը����6(��n���9H�$g/Z#YZO���Bߙī~.}�� ��h3i^���i b$�7�kW�.��3~~h�n��R�2��z���1�"wH ���{�¾Y��܀�c�CyfbF��&����-��?~��h�n�AؘB:�58�Ywmu56>�7����8���Ň���hw���e�f�)�]�HX@�x��х�T-�V[̨q{c_=5~y����(�?��,�
�I�þ����ܼ�JG�
\��P�S�(z{&�����,;�h��{;−D(U��=���X��(<�ȳ&}f������ܬ�5#��t/�\ssq)<��)N�����tQ�M�zn����w��Ķ�Y޳��6�T��|��4<'ze!�:2�1��`���4{O�X�= ��}��Tk�c�+��?���[��&DO�W�YD�̽�퍸 �/���Ig����`��:�pu�]�����W�U���Q��Ǯ��4��,d� �	砥�9G��4�x�b�H(h��&���$�^(U���F����y�$I�cPkO��S���s���m8�)�C�^*+1 %L��a�!K��EA2�3E�����p��(��2��y"��	Bp+���-�e�EK^Ș3D��cIR�y ��)��1Kԛ�dŷ׼��*��,\��Y��d�49����E	�.��J��0�����\�`  �7]h8�G�+��W;���	�0Z,�4H]�6[��f-�*�2,��ի�/I���ǆI����$D�έ�c�g�,w�^���Akm%�GrE��׊�U6����ճ�v�t������-++�������x���;������{zz8���*;m�1�<P
�a�]@��l��d����%�|Ez��+p����Zy�r}i�H_C��xK�D�(dX?Wt2(�Ea�P�� �=Cɔ6~wM\+��q@��`n��������w�)�A:߁ȇ���t?#`�}����&���]���<�ô�����Z)W7 ��mF�[yO?D�mEE�QD6��)hi�C)��f,]���;�B�%Bw�y?΃
S��Zl�sێ�@�/K����b�P��I�@U�7f�^�>ex;n�Ȕ�!cS��	4�7�B䇺;pm��Fr��d�ٻ<��3؛_!1Ts�ll��̩B�yZ���5��u/O��ڢ6�*��1��GIRbNyM8/��p����\tLAL����5�~�3�H��ԃY�����z���q�t��)�����+��4�������]���䤖F�o¤K\7�0��43錪��K� ?�B �μ��_�1�?h!�^˶�6��
��.&�����F��Y�ʖ/}o� 	��;��������0��!�()�L׻�߁@t��r��)f��&��ֆMq
�ǻ������so�̂�an(#�������	9)��n��Su�����^k�N��$��'��z�j�S�4u�g\���H��	,�0��HMB���GH9d�j�g�,���ת�3/�1�_�mk�wʼ`�C�TGLC;b����� ��{W��ug��C>��6s���x&۷�Z���ON������"/�1��κn9��%;��5��z|�>%d��XHaI)���6��Yj��������15���Q-@\��J�5X1:x�������L�FAii)����f��~��U�(�9�{��8"%N$;��ѢM:ǽ��9%$�
�3P���UR����_!ߝ"h,�s�4<�d����t����~�����%��%�|��_Q�:��D.���	��:.9v_�_Js��
TF�~�ؠv��L�P�"_D�pjV�0��|H,��Cڜ͎��z�������q���� ?�!�������k��KW8p�ox-W�֦7�{;�8d"G΄�2f��|�k_�Q�毬�o�)�$$\�fnE�ԙ��k�YW���)Z1�k�p�����ي9	�|F\��N�u��*K����ܶ��~�؇��7���h`�	W��ӑ����P�yPq�UFA�->�+C<��u'��ۈG��*V���S2&%��ɚ�NZʆ̉�s�*�����Y�U�L3�����L��_�K���l�0�=��/c�}��˘x���@��ڎ�K��{n/���ᯪ���B6H�'A,�����BA��ߔ�o��r���p���p���śY�,5vΨ��㤘8;;9	�{ �G_Yq?0SH~�t�����L���i�l-�Z��[q@��C�Y9:t�~ӽ�4��М�ן|����ʙ�����/0�u¿����I�J����5$N��p��H A,���A��ɓ6�E�����L�hЦ6��H.��h�ėH�T�arq1ryYhwL�,�"n�R�S�M&с��b8Li��QD��Ks��9�q6��SN�uB˂@��'��5�x�F���6�J,�fc��O1���K$Ss"~0mN��,��5�a4�i�&}��ᦦr.�/Ӿa��i@�g,���yBB#�4[Q(�:�CI>��:�S �G�ӡ$]����F�4�P
�5�蛿�ǉ?|��Jq^���W=�Y�8��"LJ��x���l_�5�2ב�3��z�	!+۱rX�fx����"Q�趸9��[�Z�*�P��ͨx��Ge�PX ���,F�?����3�%R��@º��Y�<#�ka�̴��Vx�V7���;���'��������zV.pA�T��[a�&�5y%�P�la?�pF-V-�����(��	Ϙ�d��e� #Bo=<�:��Gj�����W5tXSH�]m���Ts5�J���}�ރNA���#$b0!���?����g�:ʓ�<=���"7#z�`{K3:ԡ�#�=FS��� 2[5�N�4�.w̅S�q� 0��O��'o�k���:��T�/�9@������5b�n�&@�:��9r��^�:����PPۇ+t��
�y�_�@�:-���m�ZA,�;�5=��+�W)LjB��5&3�X^���w�j�:�l��
�Y-ܝ�����4I��9��-x*+I��B�q���DA��O�?%e�^��v'�a$@v/]�;,�ʯ�J�o�(0�ʃ��5�	��T�����@	ǌcw#��hR���H"W�X,�a����[��Is-�ƊȜ2���Qi�Nv�Ci�W8`�L.V�J�a��	Jvɏ��C޶����f�M�qȫ�,tf��=f��F*�E*Ѩ��������'fgC���[�$}}Eb�.^!�.`E���b�3g�����ˤe$���e��4���S���#�_��"�	[D�NGZ�.�d�Q�H�Y�%�)NNN^bW����뙦���@��H׊s ��.��e��]��!]�j�������OF�Rz��i��$���ϭx����J?�VD���Q�=���W��%� �!��!��1��-��())�t��]A&��IW��3�K�:(<�R���Q��_�_�Uv�~� ��d���Qv{��)N,�{��3Ƶ�u�Z�a���'�k�Zr�z�x+�k����?�o{Q�����Pt03BܘR^���y��cJ�i���H��s��� ?�=�oo,	�aM�oZ��K�v@X��(���e�ۊ;����tk렐Z�9x��C&oVH��#�2�Uيc{Ӌd�*�	��o��|ᠣ�z1�Z 3���>��#Fra*^WK�?+���w���� �)�S4p�vZ�۔q�᚞GԒ��Gܿ�����_�P����l�x-���=Q��	���e��Q��B� (��B�K4Ѫ���'�3��-ݳ����r��(i|��,�|f¨����������B!}���&��!��ϴ�.���	h�3�W���d�d�d��d��@Sww%���CI6�`?Ml�	�K��2�ߛ0���Ɋ�Y�X��.T��)/���eP��#<��1��2��!�W �Z�t��÷T�z��%g��bZkE�o$>7��������)_�Ǒ�+�O;�1^�tZ���[�
��N1�9U~
�B�0>�<�7Wd �'n4 l������@�4Ux�l�p>���x�H�������P�%���%|�,�5 ��Wc��+*W��>�����bF�>����}�rcK�׭w9Z0{�����H&y�7�-�V�p��pc��m�x8�jy\ޝ��w�d8��L.�s,Ч�~�@h^��4lϕ�a'LP�ճ�}sF��q�5��"�,��c6YR�z��fnja�r%=(3l��B�n�9JVe�q�)�J���m��C�ۦD���쌏��'Y����^ /���u����f]Q��-�+��1J� A��x���?财���1��d��rI���_� �ʹ\��\c��&��8䌬w�G���~���WQ�r������ ��Y-�2 >·��U�*%?���X���P�a��(�/N���&Z��Ac���Y��PEU�R���Oo��T�µ{w*$+�J~� nv�F��Ψ�+D�`�A�	�G�n�)�UQ�ht~˅9�䀋
�t��I���1K՚`�!�`'� Q$���Ϟ�#����<s�[`c�'�Op�&i�	bø��(��(~�VS�X�O��b"�0�%M�K^��ʴ��S��U�>a^_g[В�/��6��D�- ��x�l93�����PA�9l�+)>��z���`����g����[�k
�~օ��S�Cb_�����7"YPF���kcb�h��0[<P�嬉�n'��8����;�/d�c����b�z�NP��ޅ-)�r	��I0��xi����xX��r�s��>m�����ε�$�DD��"�E-J�����;�Q��D�]�6J�ha�т轎6�#������>����{���k���Ȅ{�g5�SÚK|����y�'�no/�遳&J@��*_�:���1�9�v!$_@�����!�J�d@LQ֋�w���� U�i(��r�lx�M��U��p����)�%d��V>���K� �O�;>8�TC��b��\��$��9�������7xy�c��"Q��d5��s��~�A��-N��LN�d �IR���@�NS�'��������ׅ��l���Y_� �?lB��yw�^�2'*5�(�Ց��-����ng~�`��`�p �T�� D�-�,a��"�Rs̉�IV>h��6����*�����!w�[���bx�a�����}r�{z8I�$����
 Ʒ�Va����o�����ϯ�k�䳉ט.f5��9���, !���A ��!�	Oʇ��ĸ;�x�C�h�z	m�]��5܅�G$�� �=ȁ`K�Gu$^6���S�R�Y�E�Y����Kc�����I�t5���L7"�s/�W4r�?P��3�`�qO�f �;�C�?����e�P qH�>ݤ:%���ѷJ>q-}.}�M�j&��r��[�+�-�y1��Q���O/r����L,�|?���
U�;R����q�Μ={0(i��t`t���ߐS&���&���ۍs�oO~�"�� 
A"̀��w������\^G<K�y!�\6� ���&���>8I�~L 兵"�XU�h3A��<��@U����ZV���H0\6��Fdʛ�Sz���񄫣ף�S��9'2�W�^Ú�r�ԥ��u5K_��Z&,�-��������M?�}���?m�S���Y�<%�9����vRki�g�Yw��|Ի��%'!Clxn��~�m0�A
Plp���%�˰}��D�
��oV�Q��H��ER��Ҵu��
��K����{�
�r���%$�]ox� ��\$C�P���1�,�,�R�q��@#h����O�237D�"k?> n�9�x�PXwT��¥��%�����I����~�[�3�q��6%1p~4�[��":1H�K�cL�|,5D&��T8��^G�*�ǟ߈�l���]~.�b��p d��/��w��E���2�|_e�Ȝ�V\�d�`�����g��'0	��Ck
se�j���7���,ֿ�o'*F��W�P�WHѱ̑�޸殭f��N�.�+���H�>��h�s%F�u�	��_�d��+H��?A��^ה! rZ��,�2�(�~��ǿ�3cus��o�T�Ix{��$��r���^+����p��#����呡�1J:��;�\\�H[�{��ب�z��
�ai���%<K|x����7D�㼚���Yo���#�)��U��:�>�ר�򏁐�zd5DV�#�)s��}3���+b�~Ne�35��)�������v��zg����Y��1]�k�{�)���mB5f~|���&��T���#IL�X�mH��l��OV�8bCD��3;����Gt���<�T}���{���yg{�Ckts�~��P�%o��ǎPV����	�%xG�s��NAI�i�e_R��!��4�)Y,v~<k!,��1��ah�ښ��a��ge��������)� ��d�~T �H[����WĹ�SƯ
 b,k���BDpӕh��.鋵�Zkx�C�ޚ`r!L��m����q��ǶFr��^"D[�⌸2x�%WnH~l������Y��{�\��o�J����G�ZJ��\�gɅ<~������UU�h8+.T����}�H(�� "�$�L�n������r�9��+Sׅ�`��Ef)��׭-������>%do��@�x�Fm�s�������/��vnY}�	G�R��pi�r䘂�s��{��g�����?�7�j@�<l�ueN��\w
�������uV���m��a��k�����D�K���&�i�s:�mp�m�A$�T#h����Џ�7���À/��p�&V(U�2� =F|o< uH!�IQ�����k�W�xs����A����=dD>^�,���`�P)J,�}�I�^Gۈ%��	(~Sɞ��0ᴑQCԝƀ8�p�/�tNǖ�����[Kx�:��9�Β�+���u^Ѫ��El�Lq�A��w��`��<�
�,U�8%T�c�8����ӘG�+����%�jM�L�;���t�6���3�---M�U;�u��EyMO9@��v��i�L���������,U臢c�	yI�1�T�����¼��l� R%|�4�4��һ�	R�,|��ܼ�H48��a�����DȬ��vi&���z!�_*R��~�:��H�5�I���0�aJ�	�rΩ�n����h�����y���u�\�Z�D%0�6د�US*0H:�!���4�fn�Cv�����'<�=�L�r̀6V1��uYh�����X�� ґl�Rm��B)�l���q��<���įN̨�V�����|Gl�黀zp=w�u��n��+[�^UO�uIV�U�qR��o+J��O�P��e��y��c�y�l��τ[�Ʋ a��Cϭ�=��e��z.�����ZN��GN�u�o��Nd�ʋ�Su��U\�����U���� ��^ ��ஆff�<�� ��K�UB�/bw5Oϫ�u�$KA�g	�w�TR��`6a�+}���V9r_���
��S$x�;�����ؼ8���8Ċf���$�)7DH�m������.Y6�񽧱LŖ�{�����Q�zW�Uz���0��I���ҹ����i��n�'�DT��c>GIj֓�W��'@J�k�iĉLjp�(���yo���C~�/��H)qh�bp˲���q����L�	Li��U�n�_a��F@��M$���9�"x��S�|o���iL8/���Oۉ�r&�t�L{�)ӕS�m?a�'̃��-�𰗧�Bh2A;R���k0���:����VN��g�U��B�R�+7l����V8����x�p��lf�h?�o�Xv}��B��M,Տ6h�$Wg�}+W�P�~��yˉ��vPK��G��[�����K��X�����Qp�����g����H�޵�#��a+gF�����X��jݙ�C8���ӒZ%Ͷ��;/���U�j6��9$Y�4،<xv��;S�0}�iW7Z�A�𓄈���?�KZ���7����kң��B6���z ��$S�xE�U!�3��w�8����<»l�	{��5g~���[%�����ؠt�e��G�b��&Y�+�Q	/6q���66�7v^-m��V�ӿp����n�x$��ѕ0�ל*�HT���g>�I`J$E�����un�x\�n�BK����cޮ��PH�����Z�f�v�.���=�UP��'bA�48p;?�I<5�-Nт�ͷ���j��������$kg�?�Yo
�yn�W8�g�l<�#�k�K]
jrn�)�����������bq,X*,D���ZYi���Pz�4(6��]��I
����b.���{Q���E�*��]�����+��{�/4ǡ,��>'+6)�N�S6�y,�}a܎8�v��b������ /{�8�p��$4��w�*�g�i�]�f!u�d=qi��on��wMI垝�"9���$�~vg��[�G�m3�k�#�$H��]�=>O�T�^���8r��j�T�&z�zϫa�cz��:�ƚжݧ0�9�!E�VǢ�"�Pwا�_%�KI�#���X�ٿ����r4��hߑp��5|�3(s�N�����e���[��+��dL�:�3�\�?E�����	,�J�D�Ӡ@�QK�x����WH�^x�6jإj����G�v�����E�b8N�OX�3�(�q��2��D�K_��pvRjE�d�jQ{_T�74�E�k?|�ΒG ��7��ݵ����DG��I���H�S>�+0��R$�D�����d��gg�j�ƊUh�S1��<�z +�&�����D�=�֢0�_������o��U?ܚ�D�S-���L����d�` >���/�Y�abM��p���C��c������x*}#B�~���Ձ'���\�+(t����5��������P�S#���3��(��
j�Z�D�9V������ޑx)s8m�������
�������`�7�Ӣ:�b�۲�[��{#[�i߮,i�iʬ�^_�%Я7�3 ��!��B��UoYU3�*���,�y;�Ǉ���k?��~~����{r����	��w;K�vC�����fp��Ș��E�¥�$X��)h>vb����A��E�l�ES0E�7X��˹�O#�D�����I_zH�I�7�R��MS�y����yv����B��v4-0"IZ�5{���4z��2>DN�ϯ��O�z�f�G�~�=�:>�:�F{�^}|D�sr��w�#W��)n0��Z1�E�}��@L&��4nc^7����y�<�Ȧ{��B� !�(F��H���Z��"�K�9��.7ݽx4Sg��\�`N�ϵ ������ՄƁ~g���C/��WS �X�_+ڶ���%&��ү,t�7��p��%� ��Z
�ri�~�|B*"��rP�Rq��R4j#�1f{w��W��J��~5f]C��k��r.~�3��2��z�Z��?����3�3�m�.��Ȱ���C����,T�o�#y�2��@��Iʺ�,����j�Ӡ�g(*��l�D&/<F���H�e����|(��3�;�{�gY����]���n����{v�T��~��k��հ�!�!��t�(3vA�;�>��H�s�=�q�2��a��Ej%�j�ޞ/ J�����{H�5q�r����;��X����d^�霷?�e�}	T��x펬LtZ+%�i#���0�D+ekN�e!/���EL�n��,^���4H�'�J������F�����M`��yw�Κh)tG4p����(+#*��E��J����E֭*��b"m�Fѹ����h�JzI���	4mԝ����� �>>�t��i�T�&��*��KbS`�r~����v��p�⅟kv�Y$�m��#�m�ݟlm������9{~�����R�����1ϻ�;-�̓�	�ͻ��F�,_�K��_��;�fm_�.�f�|?0���T����(/'�d��|��3� �~/,�k^���	K�����}\`~ZS\�Z�~���K�iu�~�ӏ)�%#}س�` c��@*�0�K۳�5Y��2�Kj��0th������$QV+uUuW�ũ6��)���1�r�}·~�뇤�/z�'�c�	s/~wȔ�*!@6���C��n5���O3���y�8�ծy�ó���X^^nL�
HqV�b�F@��x�jKK�!s	��'�������g�����6q3����O�|�/�d�G�ttt���(���ٍMf�&0ڣj5�j��d��ϹvO�{�i�C����Med,e���©II��Un�=���]2���nԽ�p��l��g�/Y17IF&��IePx�g QW&�;�����'�a� K�>�F/g���@��~<�Ho�?l f���G|+�$66��U�G�Z��
�9�e/�vo�ud�61�_W�<�ݭ]Q�눿PTzz��B�F��IH��P�r�Su�����t��?�F�Ww�t�U0��SB��tl�gW��+�IC���qE˹�LX5@R��A!j��{B�"ڥ{�n!$��%~Y�F!$�~��x���-mp9w��s����8��@;pQB���|S<����G&��e��avE�;�iJ�gĺ`�H��W�۳�r��ץ���I��}���ˏ	�i�� v��`YX�B_�4,���,Vg	7	W'kMp��#`�<|wiip+'ArX`_eD�ش�W�vM)G�+;J0O�}�.�`��|vDr�U6�����(Fmf�ͩi@��#�vK5{��*n܀ԑQB�L�pwo,�E��1G�f,9�[�}���)�M��4oɿ�.��O��s�w�C��K�ل�"��f��$&�s�{��*L�e.:�𘅼��7u���BS����U�Z�8x�4�Bmv�0��;ڀ���#�6�����ￆf/���7� �x�[  �t-o@�cq���U�q�d�8��]���< @u����k��n�$�_ Üs�Û��r�������+攝_���eb�k"�/�MP_.��]#������H匓��S2�����}I[[�{������T���`/��H+0ᵅ���;�S�E&;�J�5��U!�9%A3lh Z����:-&1[�T����[hH�ܜ(��^� ���y3d'ʔY���N��=�	B%n��(��!�Z9��t�m��j�$|)�/�L�7�B��źz����=%W$$����2�@�>�M$�Rd���Y$�rJu�x堖��+#�49��Fj�z��y�l��= X)���^��"���OY��%�SpBm^�o�j�������+�е��\^���E���t��W�8�fu%��=�Ԉ��S�l��l�Ŏu��2�K�%�	<y�|��I���?�q���RVh�Ӻ�+��w��2�dHh��E������\*I���S�ܒ��C�ڞv`K��t�H�H��A�E+�Zos��������S�<[����nW��t��Zp� �z}���}Q,�(ϗ ֩ۄ���(�3R�_�eOn�4�?�TQ愠�_N"x�L�Hu��J9��YH*ć}S�dp�����3�O6� ��`�p�h`p]BjY�P���t�O��xI��I��'����y���]��E�:��VNo7�2�%=qu���.��B������	a(��W�#�̊��@�Q�����(�e9ۡ�yQ��h'�@�\�`ޝ����s&ƚ�@��W7t�!��ק�r�A���]�%�nPJ���S���hK4���1�/��y3X��,�I[����Vcq�mq�Qc�ת���NVv����J�S�~�-��H���T�a�A�a�^��j̜D��Gb�\�+�����%3Ͷ˫�y����RfN�:7��#֤��9'���x���ɣ]������̸�|OiCO�,�y�h7Ck����#s��sr�$K�]~�:�_��~}��� �Rvf���g������i��l����v׹��Z�Oq��+�v޾OW%Ѽ�z���W���wL��a9�Zws�Y��W�����K���f���#Q��#��+o> c�S��)r�ۮN��pb��h&It��$���ؿ"��=:jkBK�K\�[g��z��^�&�mP�K�H�sB�d&v�<��m�v8��t(@���'S�8���L ���:��*���H�Tڒ��+-�9qp�͹�V��$=Z�I�,��|�<���t Q���p�_��J���ěK�6B� �EE�>�lki�#��kfp�V?������ߴ�)��_��u�s|*!�uj p�#���/��B�	�g��)��n�P��ig�3������������R��@'A�FGt,�@T�@Wi�	D�\�E8���hF|���x�������g�s
��F�s��ue�j�.�5ִ֞��܃��&�V����/ �J_��6�)⟬��\}G�?���8k�!���)O�@��[W�RJH����m`E����ޠL�ߊ-��	��uR�ɜ�¢����3��ka�\NB�ݿ9�ɞv[�!�D� �{�R��ǻ>�5Q�.��s���|����!�<��;�_�#��l�9���� x�	��zmd�ڨ�ċ��+|(��c�)�12��"ӗ ���%���uL4.�9@�@�>�=�O��M;�d��V�zz��k��z6��=��"���Sj�O�����Y���c;�	��J�R���OLpМȈ�- �o����5��=xo���cN�2��{��"�ӱ�p�ٚ����|y��7u��w�){S�SHvx�L�<����4I�h��)����U'�ojH�kd�?*�Y}�� �h�i�ƿ�{g�ÅM<���;�=�8� 5�!^��}�a�$L����': �%�&�S����f�u���9��C�9G/r��{H	S��^���쑩+M���Ja�/�^�yr��nOXܫ�4\�H\��ϯ�Yð�)�<���L��O��<�~���!��?�h��^D�zs����N���kt�}�9,O�";�dL��2�#jt�܋�;jXd�a!�|����sCD���M�*A��N�}�|�`���_/�"a�»�e�0����v�Bc��Tc����M$�g������WA2�ą��/�q	��)L]�P�p�J)
�e�y�^�g�^�?����ZY�f�,��i��������܆��zٳe%��������_�� �M�;)O�a��1G<�f��>I"� Eל܂��ã�g��Y�j/�S�wW�u�7�t�H����ιlT�-n8J)�?|]��}T�}/�ѥҸ�Fä��¸a"�0�˶)��9rɹ-����<>�~)�3�K��礑T\S�+�����]��"�(v�P��^#iJ"�$"30GK~2k;�5]&	����*Yu���^F�����d^T���|��H�ۧV��=oO��Q��XI`)�k:��V�G����Y6�.�Pe`�Zd�ZId�ꘅI���U���8�_RR�1"�;N����!��b�nI�{��x�=�L��������0{ִ�ɧ'=�������2V�,���?,]��0����\9�Fam��q�?ZfnP��c��CT�qY�5Zߤ=}�7�q\?n<��A/=+2��x԰^ �������}b�Lf�U���*�Bv�L);�Z�Y�5�ji�p;^�	,��N������(��C"��z9�B%z�mu���,,��\���q�>�3WqU��2�������j~2�YLQO�n�L�̆����"J����J�\6�AB85Mq:σ6Mc�J��+˜w������5��TU��،����!�������m���gfh��[D5��@N�~�1�#�ןD��o���Dw!Bs%d�s,a+�����h��@	��Eœ(���r�R�7�>�T���#��:�A*t��fr�Q�*��ścFUa�͹��)��vm���!f��̥=�ʽ�Yy�
"��\'`��NI";��~�e����v�c�0���#���Пw�~����8��,- /u�$]����؈�&�I)N�1�̪vЭ�U\ Qҗ3�(=�hկ��(d�t	���o�S5�z)�r���R�R"D=[�ۭ˽�^���3�4	I4�MÔ��y����W'���^.hfg��;���s�����k�y;�z�b�/<���'_�
 X$��wL��\d�W�y� ܤ�C�A<�^�Ɵ�s�]U�@�N/��s��5&�D���Q�J�Ә�.ȑ��:{^~������F� DeM��n-�9���r�����o%`����Y��I�9�w�|��5-�$�**�E�4?U��ib-B�����o2��-�e���<8��z�� ���7���d���K���&�Ԃ'c��b�bF�A�jA�\�M���5j�q�1=��K阨F/S��y֎Sh٠Ҫ���xǨ��Ev���f��r#���&"������i�YQD����o��W4����L��,�#�(�־)|���&!yR��9�z��x��n���co��Q��sEc�I����Nc��8N3�������)����j�n���R��8WcE��#\s����b̬}�e�b��v�Nz�.V�91m�� �qֻ�r�����WZ�<?ڲ+.��E�FbC���Q��JC���۫/�V?>+�����z���ʶ�&1���nfNm_֜����-�԰�sLm�M�SL녚�if8�vFUŵ���k�k~{*�b֖���E����� LJ.Nz*0Pf\^&�����t��ɖ�;=�M���Դc�'�8����5���YF��f�~s[���O����;'�7�53fǌD���zy��=I��ζ(��F�e�Ȏ�=��w�E_1��K���l�>`3�c��'?���1�ǯ��(�ְu6��A#��K�o'�f0aP�3�� ���f곁����0mH}h|{S��A��ݒ�[�9/�����P��G�Pr�����+�/O�o���E�{�!D��������q�
�~-M��s]p��c�N��_��9��8�������g�^-��}3��;X��˷[!
�7_nEas����]d_cs�8�-[�Q/׬����i�
�Pފ
~�,�Ҧ��iD4�4C/b�O~��R����L���I�^���e85���|�QCm���k�������,�k��J���]@.Cx6� ��72��Wrɽi���=4�m�������37�r\��4��dlf*4f�i_$�F0��VO��N��pY�m�F��H���e��*�)&�E���ٗ/��o,G�M9�T(|��YR/�5��O.J�eg�Qy��=��`�"�L*��v�[��WW�F��)}�����#��tJ��.�5f���"����	����K^�)�ń�Y�e�E[����a�vJ�4_���~]�h����"�>ן�sJ�X���.�^����s~&�b%�;
6�I c��<������%�nS.u&@�e�z����P���p�H*�45(�'���=��KґU/oU���}+ KʮpF�7�����Y����.rܦ�%�E���gL?#(Z��7�����=�6w����ȝ�\y�3D���7�~)��9z�6�^���S�Y��ձ*0#x��.w���F������Nl6�w��|�����Gis���3K��$���J�W��us�x!��L����F�f��,WGz�J{3�?�������?��6�D�%�� ��v�n��	��d,�X�~5L��Tvz=5��t7�����TE��nm/�x�vc���y��l����5?���:=b�F״��5�X*R�k�9q:\�]j�q�U���5]����T-�&<�r��ާ�!�4.IH 3|Q���\�.���]�]�#��Lc����� '����\ը�3#\�����^�P���&ڭ(A��5�/�I��jz���w{ZI�u��ȉw��I��5j�W�l��^���3 �ȑ3ӈx��:g����G���&����/�وE��D��: �:�R��M�e�FR�_�Q�7��\�����zp�H9��C�ҥ�I(-y��kg��Y3�C$�de���IL���'�C�� Z�_�N��&���XH�s�D��xD��z���a�$;��Y��������ҽ�5���䏻�Q�l��PhZͷ�iu�����Rì϶i �|�NW�T"1>����ƾS��%�#j+�Qkd��U�`�ข��t�۪��('�W����̰Im�ġ�`�U��J-��D>�l��%+��O��8zE��u����E���`l#�>�6W����fTȣ'���ʔ=�N�'Չ�� Sm�sf��]t��b��\a����T�#�2�{��Ib��)D�JZRȚh*�z�a7�BWf�x	��
+�z���r�}�A�gN��)zѺ��f�ڴ�`�FD�?V��[�\�a8\���g(��yS��--�h��26rr�������(��������Ym�ѳ*e�dv��h[��I{ɨ������\	/rŸ�z��u��'^��t���J��4,ٿx��5W�6A�:��&�*�`�[Q��4%��ڿD״{�[MT���"t�,�*�+b���A��jWP�ӕ5�!��>�H�J{�~
S�h�3Y�.F�$5T�57ؿ�gD�˭��F�5���Z�tu̎�=��$���j��E�CL�N���ᘰt��.�F0�f�g�5��>f�c���Z2;��*г�Xu�\��o[�7�q�Q�6c�œ.����K�]��_�]
�;6�Y��,j�ڕ�]���=�@��6z� �v��k�x�����3�o��nV���e�k�w�l�B�N�F(`��Ŕ�j55%̗L��<ཹ#�ͥ��H"���;ﲬ79ӯn#�J��4<g����ɰ�,�z&ŝ�-���U����Tz�&���3�x~ś�����)z�_�HC�5W����OEO�^*�z���X>��*%���Uva!⺿$��2�b )���"l0�e%��̻���7c�F�/���:{y��O��gE��>�|"��6-��L:)=��뻁^Wv�{���%+�o_���{���!5mb��h��l��bK�9��	3|�el�ky�Z��b�$BV2o	�[y��jD�(��ѻME���W?���k������˻ޛQ���D�FŠj�߱��w�/�w�0)��i�gP����=	�tK�iιH[�M$�JP%6�a����|�K�sK�\�A������H��AԬ�V�ط��O� �-?;���R��5b�ܣ�/(����T6�)ϟ�=Ғ'j�*�s��zM-�*\�?�-:�k[�{��j������3>����4X�^q5�7z��:�l���T+��3����d2\��5�B&�jW[|�Kz+\{smez�2��$��X7��KZ(�����/v[���h��l��q-��k����}�E��������`f�`N��A����\�ppWRe+HM"AC�΋e"��@Frv7w����n��f�?E��Md��3�^��^|�n��:��=���=�]�2J\Z�P2���~q ����Y�׽T�sƪD�f�!����HR�D�URۋ3BZM�4�u��c�mJ��������r.�34�)���[R�~���(ql�2 \�jGӬ�85������;kV�Fg�wJ�߷��G�f��:��^YU����i��k��tB��5֨%`ֺ(N�?�.߶v��/���-;��rev=�jp�ތK}<5�×7Q�8(%�um���[1��=�E�1E��O��_β�,~�?�!(��
��O��eS����^V}��l�-Ϥ���Q\�+&���tGj~�xn�g�� o��̟�ǓsGL�ڰ�0m���_t�&�K���,��A�gxw����N��+V�/fVx����Un�ēY��-[tDzv=�{ Y�W��}��Fbɯ-�5��I��<ǧ�"����e�����R����7�?��7�{c�E#��K�$���D�{˷�G>2�6�C�*�ij�p�-�]��Xad�C��c�?$QGY�(s<�����ˈO�'�d���X����q�U�����S|D�����8�mI:cQY��̼�BM��ب��o�g_Ҭ����-}pۛ�+���|p���*37�.�:�Ƈ���$8ު8�B��X��9�>���|�t�#*�s'�m���ճ%�Y�lr�� Ɯ��3{C�O���֩F������6�4hح{\uHW5�=R�i�����m���g%m$��~�R��s���C���~Q���
�4��n�R�G����L�	*_�."N�M-��V�s����p�U�	��;�b�J�xp
�ZUe�j�}f�/wN?��5���#+�:j�rx~�=��YU��_:$Y�)�8��*�£�@X�����1I�*>���<�w[-�jn&N|a�s�I?M�_��Y/�d�j��3SX64u�����!�燜}eM���^�U��qB&���8�x��V�����3,�Դ͉�M	b���%���xGe���^��ON�MiZͭkb�$�q4�\yFs
��N/�du��� �
8��M�L�q8�X�����zH��3���R��z��e7M�Q��3�Zj����׍���Q�@Rb#���~��ٓ��[[�OZE�³��}OϞ���G.D��kZ�<(���"ݐ,f���4 ��b3I��Em��x��2��I�D��U?m��Y<����x�nizp����*��ob6'h�'��^��I�I寊�i��=�qXX�ĠA;�U�e�\6HL�+������--ĥh��gL�^P§�fc$�S�6V!��?���(�<T���OYz	��Ϡ���t ��j,�����	]����y�)�3T���f��dJ�Ta��vH��GQK��Jn]��FL���".��(�;���׃�y��j���n4Fh�]�_Ӳ�����x����Z�ɪ�^�rv�����`:;v�q�||���˲�H�ll�<��Hnï��]7���͚9_٫P_�89���yZc��M��gԡ�l�>����B��:I��݉�'f�7W{��M��bʿ�L�ge4�G`O+߿�q�Q �����r����/o��"_p�"�&���&�4�S�>k�*��ϔ��MC���5�N0	��Y��Ь[����O�3J,�K6�n��;�������5��DT ������=S��d���p�B�Q�c�S�_��G�ElA�|���b'��e���M���'5zΉ	�&M���ZG�IG����,�ɟ����Z�G"�b~���w�)�,XO���5p���X`�%7�R����+'��VY�P��%���cSCַ'Z�8�l�;�g���!�5.�Va���Qm��<Y��<��،>C��}vA��CC{x��*� �e�� l����������Z�ʆ�	fW��(��}jEE�ZT\;GN���ݻl�
��맷� ��G�����,F1��`V��
s3�� ����s&�F��^<W��&S�$M�dw�?y����������oZ�5��n� H<�L�����G-�l�<�zU��N�ȟϝ�}�ܿ
N�h�8��� �#�K(�^�����N��Ls��D#������8���iN4�$n8E#���R���Y��Uř���U_�4�q>��_ZJ��H�r��J��i圭��iD�S͑�5FJ/֩�+%�D�O�d{�{Nώi�9&E�F�E��Rc�xn�
;1cc�	�m�i<,ad?�h@�	��r���S���Q�}��ȟ�;�����X���3/]�RVFƲ�&��^�gŶ�iw&��0ă�G�-��z��Yۭ���\�SqW�{�߄����G��L�j-�l���UL���>���N�%X\��`��;ZyF��ŌV�:�y���q��pW�?�x��u��h��`��Q.�?�����	r�`{D�^vf����*�E�Y�k7��#�!��.kˀp{����ʧL�~m���,$����ZW$�9�h(�>&N��;��6^U%٣�N���%���-�~�u�Y���$�=���� ��"�����`�'�G�C���>���f.
S��N�x��$b�(�޵�ļ��fMڣ}C�=9}:�v,�O�����ƃGO���̠�)�#�ç�f+J*�b��F�"uJԮ_	}��nj�uV#���]%�.E���@�53X�9�Z�xi����n�@�ѱ[���Qc76��9��*�@��*]\�'84�r`�K��Ց]v�~�lA|ư�־˜Ub�
E(ILnN�_s�����Ƣ����Pm��D5h�E��ޮ�V��i���M�Y���jɇ�zi�<X�w���f?����z����vc�anf�^< h6��ϰ|_�V��3�k�r�(Y�ҋ�J W��?���Eg�O���(a��
dH�#_S��
fý�"ECbHՁN�:��AVL��L#�v��p�Xw�t���֚̊b+ܣ=�31�\�����KϮ�M"�|'�h�g����Ivw�0qԩ%��G}(Z�6#�:��-�q��y0�0��O��_���{~�_��F5�6� �m�^��+Z����3\��lO�� ^��g�t�\��j�dİ��b{�N� �QB&Q�ܿ�I��lS�IP��y��	���^G�����k��D�=v]o�-�c��G[L�ݨ�A����Eb�Sv��؜�GE6���½�����y�;;g;� 4�wE�z�Xy-1-�Eu4�~(�Q��`zl�'-�
X���4��`+�)����<�+�H&�i��4�x�����Q���d^���va�Ƣ^���5ܨq��H#O�)��������#�uPb�xH}h��"g�w��H��Ѡx+�)m�� ��y���5$�l���?~y���frdDo���2^Ջ*3D�S�0 �k0����KK�'? {��Ta���"�Ǻ�"��8��ou�h�!X���+P��O@���&�[�}�;{_S\lD�l>:_��
�3>Ϳ�|r��"�8�le�1{j#0I� �4�k���M�����v ��º,�.�9j���նf;5�`���d�l �2��w����K��mYO������/T>�!�"#���Z�����I
���O^?R��;Rq	��z���mr���7[�ۀ%��?��ߺ�0�V�b��9��6�J#��pZv6�G?����C�`�3ZrPAٻ��I��$Z�#M"<w�-��f(]�����C��0!z�n^�Y��gg�Tc�h�#��E'�������Bn#���I���x4^�(��Nڻ�z[�h��^C�Wo�$X
�����T�}Yv���*t]ݽM����_J��.9*����������eVf�2NY �/<���p�}׷j9��3CӐ�N��9�ɻ�,�0����iX���O�F�ڿ����)��>팆�~f_ 	dSn�:ܪd`vXf�x�%�\!�>�B"�0�����A�R����;1�H�Q�k���cTORB�z��̷L��^nv�ަx>��5'�0u�Ā��lBW�,�
����<�m&�:Q�`��M��g��u힧L:5X=v���ƯN���a���lA���x�w@ߞ�9��:��A�"	��r�X�S�Y1ZaU��zq+4��6(��݋������fA�\�3�Y��.�ftl4��MGpQ>��>h��:�ԘV�k_���׾��C���ON��)�hEʚ]�e���e0�!���,-�P��c��+2�c����c섌e��۩��\����s]���]�羟�r��L&`NZa,���6�յ�?��N���b�����8B{�����(�}�����N�E��uog]�Vd�����%��>ĭwBw_�G���އ��UT��h�Wu���M��D�1��Mj�V���Oy��sێ�3���,�^e33�l�IT��I�|�����/<Q�N}\FOr^ttc�&�������w�Un�G%�%M�m���ѧO����+1�O��"�w񽮮�K���a��U-�+�k�����$�Z.�tT���+�ZAs�`���G1��l9KӰ�hc�W����*���>��b{��2Bi�4|��!�]�"�°���f���Õ��Ϗ��j�wP���e}㏞�P���l~���Ş�#NFM��|�zLٙ=p�Y!]��k'K���ɓ;�[��N�1{u��-������ez�ͷ���\�B�ڍw���P�>	:���n&�$�e���ЖRr�=�A� ]��?�8@+��nc�)E �{F�6�z�8�s��G7�jFt���6>�>�ؓL1Kϒ���:�aq$��������u4��e}3g����Hr�sk
H,mV��!�8)Z:���������,G�/�(Nޫ�44�3����A_�>X�o��}�����?��?{��Y��K�����Ԁ/>�rq2�@�X��s��L*�NK�)Ա{�h�^��1A�_�Aίu��+Eߝ��ɨ$�6��}��JJ�	C}�)�lS��NGEv�=٭������Ab�����H��������9Z�W���h�׮�w��S�ڟ ���RJ�5�/s��k���a�~�s�qYD@��E~���&�F���9�ۋ�-qZ��������//o4���<�ZtQ&'u�Äg{�!�lo��&X�)�LC��JR�t�;��Kn�˫���|7\�
.�`��KU����U�6
N��)���S�H<��49�*��e!�L0�_������z̾6|p�;�
S��=��I_�.���?~�]a4Nܸ(��Q�1zS=�WW���C'��"C�eS�c�F��x���m�Ff7�G�=ğ��4	�h��X��<w��w��E���kȋ���E�;��!�u�w�Q� `\�:چ뱇wo?���UY�P:�jZ`BY���O��qv�Ô�<z�#6�hY�
�ש�D�E�{�΅�0�'��ݴ�m���(��d�FT5r��+`ۿFTs�ΘY�w),r��N��tr�e`<v������@��gܯ��q�E[sJn�㈮��v���-�����=K�fcW�R��/8���^�����HE˳LLPӫ��T�F�)���
�i���%�ǈ�~J��s'�${��\�q��g�L��8�3oD��z�Z��:�Շ�o�T��"Ն�!��0�|`�x)KMIO�0��9���T1*�A?���6��hqH���s��۱�=2c��w^�t&6��⡥(�6=p����7,eufDuT5���!�F�(��������<�U�����v���&u�'���]�MC3���m��%u�-kNɌ�P���!(\=[ÅKa�����F�Y�Kg��k�J�	���.ƏE~�^�1��XS�}7�������Q6��v$Tݏ�M�#�R�����9"��G�=��3n3n����$Xd�j���j�P���/��m��Z�lы��Jǿ�|���Cg�l�z؎���?@�Է���m��y�v��\�G�[�G�}!Sz�BI�ЄL�7��#RVIԽ"�7�k�}�Y�E����f�/�?=�Շd�9��a�D�F�|T��������>��Ј�Y�5(�ittޫ�l4X���"������AO,�PVɥ��da�[^D�{,Ƣ���dW ��0��Qswxҧr3��@VYI(�gs�{T��6, ����X�ߐ��ho�	�/$���B�D�?�oįq,
k�Z�?��7��&z�E�1��۸x�*��3�wtG�����;�S�J������x�c�<[ҥ9�	�i#��<�ц�����`V�q�sU G��0�H��֖A����J�:��C�@�5����Y#Ӳ��Z,�p�-��I��;�"m���$v��2<d�7�/�>U��b{��]]ɱ������hլ�%o�����d�;��/1r���Cr��+.�Ʀ�E{��:� �9��Bw{���v��ЃR,��Z|M�6��WN��}������rk:}�z��ڼ��l����Y�������>���d��߳���5�Mj|!�@Q-P�ۡų;��5�<	-h�,K��yM8��0�@}͟� u>}�)�ME��`P���oz�-
k��:`(ix'F�߫�"""�jf��Ij"M2�B$��/��P��3�J]pC!�#���m!Mf��*g�?̍c1�\ c��!����xO�r3�.S�5��I���lRگS��.��N~F,�*��Sȷ�l�*�)��Y�l����	�L����{B��K�y��a[u=�f$�e�d�&FWt_�-�_|�X��8~Su)ㄎ�0l���B	g�����E�.\F����� C΅9������z�b�r-�RD��o��QDΥ�E��) 8E�b�J�&��69��T��~ź����KiCN��%c1G�<�F�$�ʬ_x��+v⣗\>B��z²ө�h|��� �,ƀW����3�%B/z~����]|i#U�1��)6B6`�}/�� 5����%�j�O�11$������yC����o�9�,֣Qo�hZ��@���N-�N�Jg��q� K
��:w��}b"\�9d�R錡�+߈>�R���kg��h@�|�$g�O��8M�K#J�V<��4�o'�#"�2���KFdٵ�S����L��/�ݦ>��������c�$`N��:���`�[lC�kY����Nظ�O�XMN�D��ҫn Ɣ\ܯs��A 3|]X�髎Y��,���K�&������Α9/}�'�ɭ��ʭ�Ԏ���N�`�����_�}��^/I���ƪKm�v�l�3�k�c�!�\��s�.��KЁI3�����A��2��5��vIy�Y�_�E̫�eIy?Ϥ�l�e�:�~`���b�v��Ȧ��ɵq�� �3�Uɭ�?(f��1�;���A�u�.�Mf�����Gr� s낙��smm�-t�Q����=e��S�%c�k�3���{.���������/{��=fLm��+�~1��9�2�Nc*�R�ţ��o�9� $�i,�#�rӢs����e�{��o�i��&}G�:�N;C�8�>8����G����d��c���ܿiM1-#�_I#L�&�UB��� lk���X�,t��d�D��lh	k���y]v�z�<}Ǭڛs�;CkY#\����}��gs�z=g��EM����V0�٥�Z�Kך�����.�g��x��c��^�w�q�[�*6�U]g�S�Ig���	Ȭ;C�D���?~���ml?T��9�gR���ǕX��-vQ��qU^"c4�}::��[��eɇ�D @�^���Xa�g~�
�g�����H�v�ݶ�N))���:?%��u��zdy��-QQ���`?ۻF�HC}R
=��]�����h��<*�D&wմ�U�Im�L��^'�Q!+�l���cQ���W��]�%1H�m�L�8�s�<�v��͜nk.�� ^ ��B+�-k~t*NWx�~����h��v�.�4�/a��9>UG+W��fz��F�#��˼�,�X�D��u>䜍$�o�up.��02ˠ��� ���4*�VW���k�*&M�;�_u�W��K�2j����Z�,�5Z�VKI��:��ԯ�rWCu]2h�pEs�xk�pW��4�-CyX��۴�r��`u����P�'4
Kj��I�b����`��ډ\-��U�YK+5�D�d�?'H�'�:8�.M3Jq�H���Zq�I�8�%�Ȕ��ؗ6�DӦ�W�k�Z��)c��g��Ք�$�\QΌQ|CN�cV��dZ�b�[|��sIJ;���W ���%J誌�3-��Z�Dz_3ZX�U���n4�B� ��U���`M3T�m���@��yǗ�ΰS�������¬�Ii g�30�@���9?���S�!�`}��\#J�Θ�l~U�B)A]/�3[�߿�j��bP�U0�z+���"Û��Us3��W����h9�+4�����)�*q��A�Pz�p�<p ��*$�r("������'�BѷO/�$(=����GA*�10`׸g��7�N7R���[N�V]�Z;�$277'�F	V)K&��<��_%b-���I��<�c�+qD)����~<�4h��Z/z'���/���'����C.���Q�yG�C�r��~��%)���ωP�%3i"P���!ӛ�d�����������#s�܁V�,
j��O�p��rԳ'{�q)<Ô{�rd-۾�(ֱ�y�i��H1�5
4�I�䎶X+�L*>�hue��i!^$�g���_nx�b��%:}�{��M���kO���h�0Pؘx��J4M�4���kO(n��y3�V>����=��L[]�v�j��z��H�U�Y&(�4_x��� �b�c�F�K��`Zb!�݉F&Й�l�e����|�a4��5��ajV�B�Ky]{�$ѹ����g[�Y�������x���Ӗ~�<�L��X���Zm��o�j-<��[�#;3,w�]���<�~: �v����!`,(e~�*p��R\�'��z3�>�RW7f�g+Qˋ��Q�<������6�fD�<���~\ś��%�T27�(���	.�T:A�ɞ�e*k*�Ů��Z3�TPZ����$�5�ݳ]l�gF���9~5=����V3	�ҝ�E�.� �tbR�xP�M�|��_����I��]J��r����A	�����J��Bt��^ނ��B�`j���dmm0}t��w����^A�_����q��~����sx�~w���2��q$�#�?;��� ���o�s�ƥ����H��[�/��Gp�U�x�)���H����r�>�S�4-��Nv���mE���-%�_#���5lX��~�{/������[������s�m��I��{��7�i��]�u� PK   T��Z\���� �� /   images/c99f0c6d-affa-4fa1-a395-2aad1347a31a.png�WTSk�.Dd)*M�
���w�R"  "�"��kD:�ҥt"���Tz�5%H�'�r&k�g��W��\����koy����7�HB{����|�����·�q���|+�s�̓g� ���_��'���n�O���n���Z�<==E�\-^�����I�*��@d��ڽ'^)�ً�/�ke��{-��%��Ll�k}.��p�����\�0-Y��!�Eޔ���H�ǥ�T�����~���Ύ�-�j�؎5���������܎^N![�?���Q`���,RPx���y�p����7�ӫ��?�N/U̮��>��!�G���'��3���4�g������V�yMx�t�A>^���o~�/�32y5�i��_F��dN`h���3(������d��h ����;y]����/U����EuX�sj0��_�o��X)��+�2��w:�<Ӊo�]Hf��-a�.��]�ٟ�U�b�m?^9���ih�.�ccW�V3@�5��>�t��-|K\��4�zf��/��3ci�l�\��ִ#�*y��5�M��N�Y.���W�=��qq�Rz"�)�!$g�,��ɥ�MhC��p�_�'Ի��+*�C��,�H�[��`�{ӿ�x�{}�K�T��X<���F7�و�/�R�N�=�=*�]�9�-F�_<�|U)�i�)$�|WkW�o	ڗ�\�0��d>Jj�,��q�=E��:�#��$>�ް'}u���B<J�%=��^8��lY=�J�hAUgl+��#��H-�h��Ͳ��f��/��L��j�F

.�>�,��܌�8]=m=��:֓YDHH&W?pz�t�bү+�/�C)���������V�@��Ce0��n��G��P�s�k,ww�|%�ʖ�	?��
Ck~�.�@/Y 3xu5�ya���V�fh�����H�;�Ѯ���Po����ȩ����|�~�I�������g�fM�n!�a����z��s��b~lk�t��V�f��ν�n)�J,.~�( ��L5�u�\c���H3��W�a�x�ڟ!�2}ұDR���Aʀ1�c���}��֠���W<�y��KI�����z�]a�	����5���!"B���L�y���`�p�;\�c~pH-�����������П� P?\��I�Z�`<�O��{/Y�!��c�\Py�Y̫<���K��/h'��E�,��j�Vd�Y�gd4d�یT�3�#���L���Y�`M���7:8J�5s�bѓ�>k)#:���<`D���̹ؐ�`C7��8�P��IhW�uo�;�~ڥ���t��֭��2O�f���V�
~'S��~�5�L�1f�DGmI�8<�b����c,8��9,�Dz�7�a�2����5�v�k�s.��)aP �D�iM|���Ap�5��ww�S3~Ζ~v�k��86X���>�'��X��� "���֯֏p���}�p�fDw��Z������wXz�.	����,F>s#rB�(@���
�=���T�5T�;tG��XmD����I��M��w�W����@~�~���W/���S��P�7�I�bot1����-�r�l���u5R���NzE�/r��.�s~�%�-�Z�䬸lZ��FgK�W4H��� E '�1�_5�6�nxV�s���?��膸�������V؃5��G�{ӡC���F+�5�̚8]
�����e���W�|߷�.�e�Dq��."���=��.�Æ�L�_��-� dv%0ȅS��H�R�j CͦW��X�rz��=4sd�?q�����e80�&]��u,j�=zT�܎ͳl�$J�'��g�σ�/�2��}��4����Xƴ�:�!|�k�ҷ��#7s-���@+>�0�#�.����$�mҥp��� 2�Y��cm�n���3�D%$��<. B�A���)�~H�}�¯[��0�4��}v0����aV�g�{E�^���<X؂���3�xI�+�u����n�iV�sw�	�$JpT=(���)3Ɣy{��Ù"�.=�}��A�����p�[�t��36����mfuPNX"��?����WƭHK�>{�%l��n�F��&Z�}�s2),�G��0*�'���06bS�N�n0i��&s���?�v4k{g�����D~yx���N�m:��E'֏��}J�*�3���fl~I
�4��*�g;�{�� ��v�D�#*��`q+�s���3�݁_�	1�	��q�b�75rj�L�O	u���YF&W(��h[O:¬��;�I.z"�9s�xwZ�i3c��H�Ɨ�j4���;��p&0L�o����������(���)
=����	[�Gj �iܚ�*�߭�IO��hA�̍��N{�-�[��"h���ԑ��ͯ��k ��gV�i��r&3�N�P��e�����S�.U�����yN�f����ak*����ءu�H�;��(��5���`�y<B���m��^�+SN� �z�ȍ�4�ol�H�#Q�׀�|+y�=;����]��yv-
J��� J\�DȊ�����e&	
�8�1c����J�C3��j�)���7����³=��z�ԋ�;P�pV�	K�������]Q��*�]���dNe1%�6+`�ϬA4�a�i�����/�a݁HD8�W��鈘����{5Ĩ _��In���˸(@�Ӯ^�&� ����>�N�~�!��0����L�4zx���e
�I���k�UW5@�q��;�5���	/�cbc��IY�t�zc�JKK+���䐐�����éȬQ~:y��M�������pg�obV[ݥ�v2�7�b��9%�ܛ0鰷r]��vo}ٷ>Yag������v����wy�K�^�sO+}����U�b�Tۈa8��&�7o��"�%*�7X���]!{���)�!���nqyY�8�K����g��\���,����!mѶ������̨<V�Uә�(����e�8_�f�6����SX��� +b�/?Y���+{sγWL�r�n����n�|k�A�a%�(>6�ã��
I�37,��ԯ{[��"�Y��y-z~O���iuل��.��~� �ؑ�-����nǲ�y����Q����F����0��E�Cvv&��;��	O.s�y@箒�X�94''�6?�Ι��ޱ�eTc�2���&^�|�H�^]ē������S���m4T7*[l�˙H�5�x��Q��V]}>q�{�����I� aJ#wY���ޣd�DI;���g�*��5�x(��ȨݛL@��i�G�R �5���Q]���_�t�xH�i8�ap� Ro��h��e�
)q(Q��u��/�m������}��#��������Y<('�l�L~���S�Y��M�9y'>K ����@���c����ekϕ��ݬ]����e�K��Åwq\3�cu6F�AL�2��C#강r�Ik��?�b��{$է %R/((�}Ll�D���X�,�����gwo�9$'G;�o�P��SL��/��q����>� sIp����K�Y��/z������,��TPY	-��#)�a�+{��mV3}��*�}�
��
.�W<���B��#b���Χ.��H�ₚ���}2s2�60�H���,N�{۝V+Z}���*ڬ��P���FΑ�H]�m	�1'��f�I��d���Jߩ!���Q�A5�NOd�'$,��(� U!���ȍ����g� �M���ҩ��1��(����YS#|�s�4«���L.(9�4��ټ�ߕ>���sH��y�v6*�LTC_���|FO4~lה����MN�X��^��L����[�A�7�p�Ig2�X��wr�����gO��XN ���⌉�m�e1�;C�E���JJ�J����������SKz%7R��Pr���KVi�JoF��E>mj����l�ME����ޏ��<:��P�H���#%�=qm-�V�����8%���(��i&?��?���Bff���>+��{�_��Ԁeˈ/4=(��V:{:���Œ6�AŲ�Q�1��H��.�����YrnBg��r3��֗�,�W�d�SM�� �8٫%�;�t���_��I�f~|�L	�`b�]{����S"���$�����=u�$�c��e$7G1\�r��}��GB��O2~5�  ./=HSBg� 2��A�iۗ8���;-�A�e^C��s�>�1e���uT@H��;���_����)}q2.s�,���l��֊�u~���o�屳eA!w���] (�4��WrN]WK�d�y"E�O��g����y���_�!$�r3���v$��@e��v7���+��cΗA�:�"@������()K �"_y��Ԁ*D��M�2��\��i�ہo�M}U���X7}4�phx��lB�a;c���pXE�}���=�=_��+{��v[rZX���E����τ��5 ��B
M���,���Wut��n+2R鞙�<����v''��/���,�gġ�*&L��|����n��ÕS�/>���HV�K�*��䔌JR"9ܟ�2�8E$�B��<�ہ�tf�J��?��2`#�l�>cA����z6�N����<16O"��<6���tf�o�`�m�eY�㣣m��!S�4�42���,YW������/0h��×_�).�$�jx89S�Y�:�Կx�~�n��@��0�Mf뙠�e��M��_�A�Z(A7��:#�yR�!7�i���H����5����&���=�
���x��%^y������=��1�������ö�n@7���Ь���<����jA���k�noS|TP�:�RGӔ7 d9��V.�����VX�tL���ވ���J� �9�Y8�@C�إ;��_w`��-H��t%M�|��r=?ɽ/k���<�N����&Zu����e��?$�6C��?���l��<�~C���G�����E�_���@pሇ\q����_�~��E��8ƚo��eͳW�H[-4��!�Ӟ2����6/�t\��{�[�n��wVnUB`�0֧S���a�
���׍�n��u��� ���K6��b����u��I;-�T���6�s�ax֙%+lB��kg׎]�ޫz�̕�"��������ɿ��G�FmH�g#�&�"��6��qs�F�y��I���\�����z\��2�_�p�W/g�3[#�dE\&�#	H��K�J�nu�1'�(�[����1!d���k��}�����ܾ�����b�_ .�F/� ���o���w?�qa�z�k����ҥ*��:�����������x��^�R��hIAp�������#k\T'�rF��ي1�;$D�M7k+?��y-zӛo t+���Tf�ӯp݉�L��	8��s�̫��N&~W�7I�[Uq�<���ݝ�@'CNؚ����pߣ�e��onw9,��KonՕ�T֌�J�H�DD���ڕ��S[O�ipd�P��O�^ݏ��Md����&`� �)s��9ɝ@�s�҂5o�<g�V9{{��&�tׇr�z�b�?RJ��j�B�A��`��ە���-� ��$	�獪�^k���+QRbV������V^)p�k��w�a8.��������6��/��li�$:n ��ʉ�� P��	�<����[�T�.����~orL�����_�\���Y��I�4���^��Ky��0����*��ۇM�í8� d��6á��鲱$�?�񵏥�1&�L ����\_V����Gx}t��k��(�J��6�S��t�a��Y:���:�S�iA��"�1�3���lD̸k}
H~����I�=m�3������"aO ��.�=~�e��,�'�JX:�G��E�x�r����Z�d����=�G�rr�����d0;9O^�T./3]Ҷ�Q�<e3S�:'��e�nE��}s�������F�ӹؘCf��(�Փ����{\���y�K8�(ݶ��:�_8H|Q0�l�㝙¾_��'q�h����M��X'	�'I?�8���J�J���lD��.���p��B�����zm9u���(Z�d�U�Ո&Z�D�DQ�z�K�VVV��$ 6�T���GDEA�

��f�����氹T�Z��H�߉��R��T`�\��[��C�&�B��f�&��2ݼ�J�= a��]t���'��kkߓ��Jm|������&��L�e?-9�_�V�S��qloܽ�?[o��R{��-�:��Ӻ�^(��h���Z槰��w����S�P�������rK@*؋�f��푳�ʕ.���6 ��6�n"[66�+�P��̓S>�r�����
��%�{Dfi�z��N�����E�Ч�������4T��[Υt+���o��	�| �D��l��Ü��'M6������ d;���sW��N�{W����\�)��D�<'���O��"�g�o������ѿ���@���Z�R��fih)���:��ñ_�O���D4F�1L�z�1#K�J�J�*eE[����a+\���p�a�j���z��j۠�#��� �OZj�ۮ�1��� �H����aE5����>�� �.vn�B_�M��b-�rT!i{�c�.[���-�=�U �719�簱���0q2�ZF�V�rV���J����/KU�&��0�^���k�}Д�jǎb�9���]�je��5���,~|�n*(�Y�.~�%�s+�>��?^�Gg&������;r�䭉��L�K�yqr����O���39�D� )������DT�W��I��7oo<'�#��79��CGPE]�`i+���r���%E@�2;���w��U�R4ꥷ{i}p�A�9�3�JG����_�\B� +P��0�T&>����O��T�%,�GB�z��z'�=&-�בq��+%1����I���O0�Ԋ��M�c��E�_�E�0M�Gҫ��^�TQ����ts(SJ���F%|�Zs�C$v����Ƚ)D�'պ�cJk��(DY��8`~
��X�<�u��=�4sw��0����On��wOB�]�=��d�Bx�g�V��;��
��ϯ�&�m�����q���>�dڋ�����)t�,�S̶������s<�ׇ�cY����Ѱ�C�����t��1Mqk��o&�96@!�5���K��S��[��g��}��N=��^��DĦ���F��	0�f��?(���`�Đ)}Gx_����o���8 (b6��u�(�),�� ���Ͻ_��{�TJ�e��F��ݩ]�.4����`�����u���ete8'��/�h� G3��6Y
Х�o�X��:dJ-��D�RGg���鸝`;��Z��[=M�3#���
�em���|��J��(%8i6�ˣQq�yt�X���U�F胢�
f���u�jE��e�
��fM��rt/.���j����??��I䄇m��6�*����e�'�)=/RpZ��Bޚ���J��5aѳ����/�^����� �<�-u�P���㌬2lj���������q�#!�X3y-��8����͏f�cB�ү������CM�xz�p�Y���ҡ��u�XK��4�~�l����H�
�o�o!���Q��TD.ípē�Cx��k��AX�C�. +[�eGť+W��q֫����X�s�A�E�Ih_���A`4��gJ�3����~;)Ki��W���ק��?��;;���N�HHg#l&���"�MO��gҎ�AS�㭟��c}�{��W	�Ls�H�G��W��^��:ч��u�&��WRE>�IQ~1�����i��k�u�?@�*{m��+����Y�T��_����g�n���Z�����̥����� Y�B�t�u�W3��q�7��W���sHxZao��K��
Vu�_��Ԁ��D��6�zv� �q�F
j�Pᓩ�m���rhN�j��~��[rC'�J(2��z��U�N����^�Xy|��E�$�D�T[��G�Hs���ܲyh�Ƿ���q�ZGS���^9o��Q��/�*����Z1P����"ѱrim*4��2D;k��i�8d[uv�gejwز5��r�����V5H9Dպ����*��oD P�>�j>op��,��I|}H�z��X���h��i�v�j��dQ(��j����̚(��o��i�)�������qNN���ŉ-J��v�L�%��!�߇�C:��s�xOF0���0�@�3��]G��Q�
z��
g������1���)��r�@�+4�\IP�v�~�}���r��l6���]�Zԝ�����7Z�v���<w5�����'<������Z������MTn[B��*P~������* �[��u��M�[���T�8�����]�u����%(�= ¤��l#��gf[Qa1��\Y�����Qg��)������[vr���A}<׬��:Z��B����B:�l�m���q>�ʔǷzo���	�?긌�:��:�'$ȗ�!�u_�8c�W��n�1T���(�r��F�^��>�}�Ӵѽ{F�6Խ���*�,��W�4�5{�|廽5�T@����$�G��o�O2S`��W�܂=M����+5��|
(�H�$۰�{(�-I!�ٔ�95`����O�+u�h%Φ㋾�����δ���M� >{t�6WP���q6_��� ����4/fEg��Jm�p}��85�r���q���o$"m8t��6:.S��h�}ʾo�\�颍�ռ�d�r� 5H垏"�盺���������猎���tC���ƕ�b��ْ���[��n��Ur����qL����"��7�rwGTbl\�0�ZR�3�!��w(���������e>���m�ҽ�Kx|���|8;4�F�0�����&))��9�ztE|�E�R|$�"�1���H��W���^O���wWh�x!���z���.%���_=@��n_v��%��L�N]]��U+q�����y����Db;}��sl9yJ;� gq)���$��s�B��Z/�t2SsS�_��`	�v���7��+��Z���~}G\{};�#���6������;%��o���|2A_�|M��E�_)�Ԋr琲~y��E��5B�sy�"�ٹ�pV-��I�G�P1���������#�v�z���,�7sLo��!�L;��P!����~7���T�-4��-����q:�w|Q~8,.�%c��H����H���u����ř��%���ϥz�.�@��Kd7��O(R2 y�Nã��%%�g�3�vfWgECzL��nB��ʩo��\�T$�t�KW�r�A;�<:^������$�~?N!�s�K@��W����Nk�ZN������0�.�� �d{�2F1	���[������7�3��Y7�5��t	���f�Jը�=���� z��#%�#������g�����"y�Jv��Q����U�i_PE�_!�ˤ) ?��k;X�A�����H5��56������؝O�b��~nE`�(#�XN�iIk�Y�yb�hJ ���le����'��G:U�d�rR�b�����Y� ��l�e��K�1�@���4����[µǥV����Z2��Xߐw��;�B�?�S�>�K[w�=�"� 7�|���~|~�+G���"�ʠ��q�s�hti�D��h�}<������\uf%V s���%]j�f���H�za~-���y*�Y5�Bn�;�8��s66v�)�[K�Z��]f��p��-�ʪ*��:li�<PM>��yLq�Z��'r���f���H�=�4�C%[dP1��J�QҘ#Z�l_��(��R-��M�|G6j��i��y=_�h0W�q�.)i�]f�z:x�heia��Vwn����?A�sl�:c�Rj���M�~�@��=�����d M�&c��k'�B*�P�-�$dR��8p���ۦ�r�}� ����L����(_�f���gq��a���o�r�ɩ��wY����� ��ΐ�2]�n���ӡt��nd�1n |�g���J�#��&7�B
<�$2��u�Z�c�6#G>�9y8D��U�l��e���kl�5�]Ё�����I��<vie-��+I�H��2�t�b�HX���z̽5D�6:=��i����/�e�خ��zɱͼ������;�B)�<s3w�dE[R�q����_�&����$�|4Z��_����(2?���Cy���T�e�P��ڦ٥��AF�%�p����=�<b^��wa����'`���VsB>�j㖭�5�~�z�>�x*�
��xNc�j�^�ft����
��&���/�j3o�*����5�BK&�]:?२�<��T�u��#[4��D8s�D��7�qI3�¯�R/w��>�XQ���׈�-2%6;��g���7�w�2|�����@����ՎF2�4��lE�)�GBFkFK�˜��P)WXB�r?gL��6�E5ޡ?����oU���
Uצ2gדG~9@.��y�s2R[;X�1p:�l)�,&P�+x�V/+��V���s稀4;�7 E��nn�21��|�'�����!x|�x/++?�3�~\�3�o��If���8n� �~�YzI쎕�ʊ�r��o+7@�(���9�Б���Rw���_ԅp/����%�b�&�s�?Z����>�<t�i���S9�TW��m�-g���f��������a��H]YSRh#j��lֶ�%(�Ç TZoL�C}yJH�H�X-*�7�^@*R_e�%bv��Q��g����]�A�a�z"�o&a��^�����*O�~�l�xm�B�U��ʰ���Å���`+���t/>�7��{Ȼv�؀�~&�f${/���&���9�|qL_���`,��|���x��C/�̪U�M*7�0�I�d�Z�M��&�×=+�T�o��Ƌ�~�w,���@�7�T����L˅��������Zч�ˠ�K㷧HF��F�k�A,sC�X�N`�B���j�D�I�4_+SE�Z�F�(3y��f!�ð�91�3<|���[��Lk��s�x�*���N~n븇OmB���wr��?�]�b(%\�q(��5��=�!&'�����=�ɍ�w]�ña=���%�Y_D(O,���w�W��4�lLC3B�{�����Y��X��^���|����ZT�E����TG��Ec1�P<���B� �e��_	�&��~udJgEjs��O���w6��JϊO�
�#�n]�	�r�G@٬�F�0��I���o����+9>	]���Eu�$F��q��i��(^zf``�{8�n�?���R�����a�cD�l����ؿw��ςv��F���#i�i����הn�8��u�dkLu���m��M�-�*,��2���x':��6����t��c_�v����ǜ��z��6�3���"3�]���ύ�j0�{���۹�H?t�Dn�0���8==��4	�Ќ��HqO��H+�~:'�7/�_WT��+��
H�dT�����ӥx�V�q�]�Aê��7x�#�QeNi��<�9%\^�d�M��ݔ��I������M�5/	��i�LNv�A���4���͐��:�i%�q� ����{
��|�|LH�������G�#�ʡ�Q����(��{�CW
_;li�[�?���Zsؽ�4��f���s[
�!�*�{޵��e�C������*9�㿽V�p��n)Th�Su�\N���wu�>�6@�bX�>VG�KtH��"e�4k�~
OR:�`I���/vW���X"��g�E��|oΩ�=����w�+����'.�N���;�i@/�u5��z��QS�,Ԝ�<��μ���7�>"����KyJ�ֈ����ԘjΙe3����I7`��,P&������3_R�*�����5�q���)�~�W+����eaoh#	�5ys���9����e�Ҝ?�X�9J�;���m�0<����Ʌ��2��}J��U�u�4���%�
��:hBǸF���utO��j�O���R܏]І�mS��z�29+_�p)��:��x���K�:cIj�SZ�ɛ'���Fm��;Z٭�%�SUx�~�+f���g�U����)~�(zNW<�8v��UT��ȋf;|ڋN?'�B�N??/oM�������6N�0+F��+k����5����\�On�|U�l�k���qc���m��?�bik����.Lƭ7O��Js���qh�M�����c_�'�{��,y������+?B�d�A=7����;A�����KN�D��%�[�V��1٘+hFL�Fw,s��s*�J2���i�4�K�ش�d��7�t����1�ADX�'}�G�JB�L�ZW�S��I���Ѻ�@��w��'�-�nmH��ty�e�0靱� V�u�~_���=��K�$�������OɎhb�N�6�t��~Y��͋}�;�r.�oC��.&N�Im����"�JRji���3��*��q���v(c{�2�=��B�t]�A �_R��ׇ���f�K�΁V��#y�����z��=��\ ����B�#g����=�?(J�ns���67�~z@w�d8��N`{�P��}�5+������/�tv��8���m��m��%��AUia��ib�\��9��439̒Q��x����\��E@��M�c����,JЊ�����I���+�gΑ���x߻)�w"�l��/٠�J�A�K&��z��}�I��u|�$[������Q�0��^��v"*�m�d��ZF�T�ɫ�H@Ⱦ~_���g�M�,����2���9p�=7�ٜ�k�0*�$
h���Z,80��q5��H�z)�᚟�vn�����MHO-�;(ܚ�k|����O[:�l����Eax.%�cl�����ʝD��y�$�<��L��kv*�Ϲ��D���Z5E
��lY����.�	��=ґ�d l�ߴ~����^��A.[7�
He�[,j�9��ME����TN�p�6J������yv�����B��Dc7�zʏ�I��8�i3�����[ǻx����-��)�¤`��Wʏm��#�_U=�im)��71��'�e�rt�{��❜%~��e9d!m�_ZK�$0��Ƿ�xlrrp���E����1a5���u�*�W��̦ �P�������tj�I�^	*���*͇�J���c;�54Ȇ\�����mU����1�����^ή�"?�S-z͚�F9�p���e�������ttt\�ieZ����X���i��Wݨ��yk�w�Q�ʹ.�Ğ��3Ӿ�R5���vʁ�fHx�e~���3ĨvJz�R�A�mO���Ɔ������~�)�������%��;�@i�^#���U������1a-t� v*�^s	��215�o�GGG�f��C��<*����Љ�%)���[� ���\VV�ԇ�ϙ�N�uZl���5w�q�.�nJ�O�w�܀?`�z�x}��Aup�����n�eE��wpswp�&�A��Y���p�L�Ơ�q��+߬��j�gV����$IO��n��_,����_"���^�3�Z7����2�
�e+��3Vn�'��ڳ�q��	�?�=�7�+�g:ٔ�p(C�8�mt��K��M����vx'����j�`��3_�;�����c��z���itx]� &�K���n��
���pv���.�Q�~0&��%���[.+�7ʹ
��]��o~���Mӌ������ɢ2ز�S^qa�dtp�����!���,��n���z+(/��x5�4L?G��Zh��Ǻ��"�C	9q+���i�<f>�Q��f>�I9�8L��(L7��3��gܦ�-���� 	���������g�8�V;D�P�Q��s:�T��@맧�T��.^�������n��!�Q.W�������q�4�<�>�E@	��г$$�t�!B�}���&i��Ә�ҳ۾�Î�]P2� �n���Y&Kf���T��+]۱2��>�R��Vəo��(�5Kx,^�K[��b�	S�fj��ܧ�W���]���!L&�M�TG%+ZW��Y?�띄>hp�w��u�c�� %��{�
k�e>���_L^�����w��Ά��B�1��"t1���+���/��������H�H�$�N�*� ��.�ԅn�R
�u��R��s�YI�-E�C[�ۏT�;/s2I�7Ȁ�g�8�8�O�k
���@\�x������0B}E.�{��+ȾQ0�7G��������u!�>�w�p��7ܸ��_��dVܨ3|��9���X1�o'��l<��!Y2��&N��YJ�����(�7�Y\fL�גI��G��A��5��&=��OQ��N_+���p{���:_� v��Њ���4��P��1?���W��A����K�l�I��B���1��Kt�/�������Tl4�w��p�g��mk3P��ǆb��8IϚ�L(rF��j�a����}P*JP���ة�}�r)T�柱H�ا���"��}eO���/T������m�T�e�g��+�ԭ��@>q0A�$ʀ����}�c��:��"���J}�g��4���.��������PS��r�F������^~���at��'�b�zjÏX���g?I:��@Jz��4����iC��.�9��U������[)�&�T���@��&L����㺱>3�:���<#ʞ=+����]���k@��H�	���V��+�l��@��������F条S�\��g䄤�Fnk�Zj�yݹ���BG;��� x��	?@@�͖\�[��{<Ҫ�E�!3F�р|�O������N�c�Წq��0F�XP2���-O~c$�9�<h�����0�4��*�ڙ�Ez���_D��}M�`�m|o���{ʧ1&���z����܏]����P��v�N��2���+%���?M�������M��3�q!���K,<�O@��3���n�_�ªp����]�Ȳ����eU�hDE���O�c{}y!��0�i��5�N\'�ojL�S�r�F�'�	�P7���ǯ�n5x��_����_e�f�?��<Nj�؎�>6�����S�t�I^
�C��$� "n'��N�C�٤e��F���@�r|�?}sLτU�7�/�n_gP��y���RL�'}X�%_�P�5����s*�U6�.C�y5���k`��i��v0#~�� J��=c�$��#��T�ХR�W�����>1E���z^�'oFX�V���̤�Fөp��Ї���^ d	��l�J�)�++Y�w��	�'He���b���+���~�=;����Λqu�%e4ke�UC�\��̄� el���+c�1_�q���ӛ�d�7I��@^�F��tŭs���V���ݤ�}@to^;m8���f�L�
x\��F���|�|��*�1<̱�GK��>��1��|�g^�z)(F��E��d.Dhg2-���Qm_s�1��h|�E�O����煳�;J<�x.(��1��T~��0t�R6b=�rJ��´�,ɾ����o�>13�o�n�(���}��_�+L��cҳ����Ԍh�\P���)hFi��U/���� {R�<�UwD)v�T��a�d>���@��lD23mϾ{4��ڡ����|�뭅t�\{e��W;�6.n�xz&>
͵��PR�x��m��[j� �w�Q�^�<�]ڄ���(yΖ��|���4M-\+������g��Y}���Pr���&OW��Y���+}|���?�s��ٱ4�?�I�������hH�q�Dw��@�Ƽ}��&z��& a$�~����x�f�ȴ"fa;G��VQ����/�.z��#|�7��� �.�:_^����,��y"@��k� f����|���d��i�{��Z\}:}���~�y��MH���%�fϽ�1J�p^�����̌��ڗ0t�+7%��1�Z�y�z�&g[�m�����X-��l'�X�jQ'\��Y���c�| �_�ۚ�ʼ�Q��h�7�_�S*�l�����Q�\
|�s��m�U

��3>*&-Ё����e�蔥e���'1� �����ziuxt��Zˢ�������+�΁2�����'5@��(�c�Wo�3��a�j,G�Y9oȄ��P�2�򧒄�SID��p������SK� �3���<�J���&�tP��W��pbtF'S��	�Wcq���Z���:Y���#�vG���l�P��N���ۗ<�	ڳJ�y5$��i�$�"]��#Z�����@�hn����:��X�@;�>�sׯ���D"Ö���`�w�Յ�Z*�R5^�VH)7�Æ�-�5.�.��+�ݛt>YrTc��Ǖ'��	�j��a���Fr������Wow���g�k�V �ASە	��WL��bq2e�#�J�����N���J�x���Sj�Ŗ���!q��O�֥�K�"��2�I|�����޺�P5���p����pHO^0`�<ۄ�It	L �Z_e��.υ:��V�Z�Znf�Μ���S�f�19����*=`R|M�Mp�.+��N�y�7�������)�g@������9�l軤��BL3W��箿�&�Hꤰ���,n	�Ђ�Rx����9%H��NMM�mT��w�BY{ş�±J���f(��K�L(3�Ok��2R�J�@���[���=�_�T<=_I�@�'��'��v �m��[�����nA	�	E�n��OY~��1�֛�5@�s5FZ� zx���6Q���(����'ҟ�Lxa��D��3�� o��11'hk+{���{Dz���j(�Ta5l��3Yic��K�W��M��ۊY ��YX�͠�v�����gD�#���}v�~@�$���:��.Y�SO6�h6_"�����z�2�+{��$Ç��>��ة*��T�]?.PY��w�A5h7����0��{^oE�5.~���*�q����������;�������H�� �(��nD�H�Q齆 !�"� �T�H����#�k�-��K"%	 ����Ͻx��||LffϬ��ZsNf��C��H�$�;�?RLKΧ���A="�E<}��Y��AnZHwiN���Z6}�����մ���_�F�τ4��5�~=K{5�az����1U���Z����� �W���DR�����cW���Ѻ��?�}��z�^O��a�������&��9�}V^ЁB�f� ��L�|���X>��Br����ۺlL�F1�0����1�,�������~���"����{NQu�_R`�e�Dg%WS�Jr�m�J���߽V�� x��"��͛�,VE[}��w�z|��S��ȑݥ轷���N�[�+���n��t�4�O������)<�ش>8���k�h�c���կ�3t��1�޷�+"f!՗ט@o��v<���*#D��߈�_�!�(��z�G�a�5V~98��t��=&�Y�<Y�9)	����#�A�'N�MG����P'��}eV½`נ&�܉��A�*�
��?�R�� ������)�:S,��H�I�+��_��d�l(v�c�������S�3������.@a�,~��{���14q ˘8��9�ATT���+(���}@H��˟���L�ɲs�li �==�
З�1��U���>Nฯ����pj���O�yv><�;���uf&p�6�"�S�ޜ�����v,Ip?�7����N|U%Ń���P3�Vvk�����6C�1�oEa�r$�`W�=������׏�K���떄+�(kT� �N�M1n�ku��ᑪ��U8�ju�6p��TR��@��Y�9Z����I{܆���T*����1p�yڝ��?w�j�.��ė�u�;�S|Y۞��Y$Ո�BM�]|=<
�?ix�ЌTuc0uyϯ����@����0|S����;|������Ʉ��3@S(4u��r��}3�Y��Ȧ��W�f���`���_�޼��]0G�-�_� ���z����i��>��Ʃ �Ke-����c'�콻������^Ǟj�?ۡu���0Z}&�����xx=x��5u�*�W��E��d����i�|�Na7B��ˠo���`M���9&
ܵǏ�Щ�դ�]E��R����N~Xєe��t�9��>z��5�H=p�a��=�$�E�ܪ��H�3��Q�i�@��G�f�+0�� ?�15�y�hv/#NͅdX�S�n�@�t�n��c��mm�����g���J�v1�D�c.:����,S+�?�k��/�б�ǭ��2?��}�������w�	E4�
���ki�CմUF���P�H���,8[4v�)���Zޣ��aR'�ףg��� �"ǧ��ڷ7��{t�����wm�<�A�?�9�϶�?X_wU����We$����hB�~����-/�w��n�N�2�]��ar3�D�L;���5�c�f�N\�Wƞs\���<�(!X���^о=ꋴ����hȒ{����uG'��jtGlK�eJ��������R�)JǏ����t���'�3�#w&����]�mդ����t&K+�"�_�=�����q*�Ë
���aR��h����C<O#���]��E$&t���6��}{�$��$\a�O"�3Ѯ�W��G
�Zt�hY�/png��@
eEs�Z�o=>C��$#�*P`jꑰ�R�a�����dq��E��W������}��E��aJDD��<�(��s���y ����j��sB_{���|����aѱT�R��d������bF-/���O: m�$�`���Fl�6�/��f�W¿�|۸��q�h�V�#u$�������!%nv5>���cr��0�1e4��=�>�*Fc�����[���hēo�8��ϩ-g+.[� ?�����c3�UW�7g�#��s({��3��|�fiڽ6zt�HĐ�E�r0�˟oŶ,t�q�\��<;F�����5�����76½o��jn��#�Ek/����J��>�'��m�A8���c�j�m*��Kr���3�q����-ԗKJ�e���"J�7Wn��ѹﺰ��|,�d
���R^^I�[��uM�ӊ��9�ᦱfAe��h1ڰ�w9���_\�4)���ӗ�d�C�L�.�Pg�=Ioh�l�h�?j���`�񐃲�{�����5��I*�
����rl?�V;�WLuW�Yr�SU���6P�V޿��T����2e�� ���i�ؖ���)��&�����(�����]pwSm�<�uV�ZϿKX���z8fXoW�}:��jj�}�༴#��<VW�
�uh꣩��[�®���%������Y�v/��m<6%T�vy����.�&ɦ_ˁu�Q^�x����t^�f����с���}�#����D�T�h{2FG�0?�9Z=���gs�1*��osn�:�b͉�'u�»�6�)ѴH�8��v������YX����r��_D��j ؝��!l~8X����N��Hmј��~��P�x^�U��-�
Ccy�b��t>�����~�����7�3j�е w�1ZLz}���p!��n�{�+�X�OnXR6NGg�>�S7R�5�r�xc�1�oL�l\��[t�Quw�༠}l:W���	+� ��
-'��k@�&�k7I����C�Zk Q����R�ի[����F���;%Đ�p%2�̥eTQ�5�1�LĂt媲Rʪ�5����`�L�m�� ��v�O��Nj�����0��R�v��כr�n���j�I�,O�L�K�1��C�M4N�?gߍ6迀����&�>�֨!.�m|�t��J.wZ���������(��`7�_�r~�]��IxQ��O2
��v@_��Ψ�j�}���,U�hӃ�&:Wt�8���}7��\�{i:Z�	04=mf�l�qo��_U��l�S9�Z.Xͷ�&�M���z�����$dX�TyX�ݒ�x�S����˧�	�uĴٙj�zp�s@��I�8!Uc�o���af�*V��\�� 1V[(a��ֲ���7�9���A�3L�n� M���x_��1Ƭ�O�r]+����a��vv�Z��YD�G�g����C��^E�V�^0���к�ɭ��c�ྶh���b�X�=[��g&��HwJZ�~oΌ D��UTwpU�Ru��Օr�K�9�j��-�#Ō]��H��ķu�cQ$��5!�=���̨w�]��٭ݍ�iߚ�)�;)�Mr ��wp���!o��R��+�^�@���rW���_�ԼKEU��3q��ӿ"A��7�IΒ���D�3Px�A����	�v�C&�K)P��О�}FNl4�*�u�;	�O�W�c�+��*�T���)�gbݶK������*pi�ݐ�&��h���߫�����$�OE�1M�p3���	�� W��Ms�NztKn�;�]�@�ү��DƸ�J 9��a$C�&�{���2T��=q/+f���kׄ��e}��E'9b�ҺW�?/�	���ʕ[e��0:�a����cW.���e�e�w܇�M����P���F34�}�wI/)�^OA��z{�e�>y;���:)(�B\��gGAn�/�QYu����"ӥ���T��讝�Y�����ȍJR�P��B
�ᆠ�sg�������g{'Y���7�R΁�h[��y�;�5$�������n��,��L����孤�1��<6����H����ݎ$��}�U�[��*t�%�C��p�y�z�ey�� ��$�>R���ԋ����ҿe�CU�d2n-�3����&ن��5����9^�D� �*��bߖrڰr_A=p�
�%OF�&�ز9YrӲ�Vv���m�2]QTe�j�%w}+��`v��rP�B�_�˷�7��002�d��^Q���E6Дo�k/kz������q��CM��<h1��3nOr �/�x�$�C�\K��)HSϹ����aJ��D(>�6���[LQ��9���bUmwy��0v�:~p��pƤچ���T���/��Uo:�έ���O��8Dn��fm�
����>"k��,���[���/�2H�b�]�d�t^�,����~��s�Xm������&�`)�nNrҔi�X�o[2§(W?=>	J=o���JO�}� _{u'�v��?�h�ФLi^'T����u��x㻝�$�<���x���r3toɛex��2V�vթ���z&q74H��0�f�̹vX^IZ|;w9���b�2b��=���%�VռD��`��BX Z;)7��2]F��Xrg�R>�}� �[�3��av�r��L�z��`&�z��S�sRb�'�,�����W@��u��v»U��ِ���n�â�1�k�F;K78aI�4�)����}��Z�8(��X'j&������|2h�I���	)�,)z���	)��0e#߉���貮�!>�v�Ҥ�������1����H���6j�ˮ��;�7*��V��c��)6���߫#���D'�����s�Dym��\^�#M���$â��N��I�������3��ޫ,P��WbH1����XXǙG$�s8��p��+�e��j�����\�?e��`�����jQ��h,r'+n=�bh��9z���HT�wA;�y޲�V7>�`"D+u��p�ø�=�Llcx���gT�:pq1��M�l��e�;�/�G/:�rQ�yv~�|�Լ�eD��&��E�&X�	�_�0խh� �<���k@�� ���[�l_�w�I/��ߵ��L�0�� k����ؑ? ���������l#�/Q�4�v�����w�&�Q�z;���#/�� d�d����S����Ř�nu������c�m��qm�L���h��z��Ƙ�5��k�h}cBW5l�͐1��y	�Q),�d:��ۛ���#������ϭf�*�|յ�=�|}�"���x-�Nٔ��G9Q�m�H���х�+4��l�(߯��c�D����%�mf�u�qP��b�t��t��?=,��-l	������<V�}|>��Z�Q��
��2�+	^|㇌b���WT�]<"��+����C�f�xق�5K!�[|��M%ݶr
�4�G�?]�|�8��	�]�[m���Y����2	e!�>w�P���|����U]~�!	 V�?��K8��G���G��>�a�UF�ά����M��1\���.%8,;�+����F�4�61b{n��w�[Ղ��,������>�7-*�^o�ZJd��b�/BQ���ދm]���� P+��jQ��fQvt����8��զW,�>��7��]j��5HSɅ�� ������^Y���a��ag���D���!�Vy���~�-WW���p�B����e�j����v�%J�׈w޻SG���VD��|��~ӽ�`�1f^�i����ջ�G��s��(:�D��+Nc}�$���/�2a߯j��bh����/�?�u`۶6ڑF��VfC�Vc�o;�@�ϊQ1"����(�%XeH��m�Ce�k�����3��ƻ�W�� S~��e�/��ܝ��؛�m垬�ծ!�c�&�L�>�d*x$�.g�ޖ�� ,��z�d3�Y�Z]L���&��[�4>����𹐴��t9I\��'�;$�m˺�M,��R'm���S��9h29FF�[߀~�]Grd;�����r�����=	��ּ��j���Z=�yP�`��^c�U�X�wЁ��ov%/�xOw�o4�,"$�G���e\����M[�
����!�}wG���NgoD��5�CzB�EebR�E�߽<�B��Qjo�-�����2����Er(���w�(��"/30s_�^@��=f�����5Ŏ�j�B#-?bVk(i�g�>�t�'"h^��zrD�ma���y{�p�
���XSy.=E���/X���Uiy��Av���q�-B\��S�nU�5 S�W�i&�:�E�G�79�L���L���·Kpұ\F��m�;ڑ��3�(��ˑ[Ȣ�ڱm��k�3���ȼ��^QY�#y*�}^H��*�9�7�F?K�_u��j�i�L*ׁ��gM��B�* �ڨ.�mE�%�I�*,��
t��8�gS��D}���K���I��o�6��^���/� %��i@��6�׽�7#k����B�g���8E��"�ca$��;W����Z18�{����
h�h<��3����S���T#�-����U��[扞8d���:�Ͱ�|@.��Q��������~����Z�^��j�Ul+3Vﾓ�>bh:_>�E���n���X���6�w3ra����6��B�����!b�ل�>1VGGv�����j,`q�.+T<���)�(8��C�{�L� �xdgw{�7fM��|:^{��'lz{t����hxݞC(;:۫��h:;Ɏr,k.��5S�*ܻ��[��fq@c-�Q�uc���\��I�dq��p�I�����G��TR�3Ɵ)�(�VrI$�0���z߉ph}�ɹ�߁�Ż&%Bɣ���W�������e�R�Q���+�h�{�O>2�VB��XTgG#A{o�Y{'�~���r�k�,/~��[d�#9Z2Lh���,}9	���3�;�΄��~����|��*���1�i^�����:I�w�^�����,�����Ę#[����E��j���t2@>��U�,G��? ���R��:�蠋o��������I *r�f��ķ�>�0�|����j�,Xe`آ�(�#hH�j嵇�mc"ģ�L<pߞ��O�>�X�Y�\7(>�&d�y�w"��<�		�?�j��M� ��0k�{m LV,���dp�J�ݕ��Ɂb��k�.ϣ�%Hp�:]j��f��E]u����S��ԛ�{~��{��ՄƄ��l.�޷f�;$�T_��iw�%�s�ڙϒ��~Oş�S�>hkk<fcmSVV[��ν�%���8i?���E��I��/��:Tg��A�6ڌ+Nɢ{�nχ�J'iA&%�TA_4G�ʔJ%=�p��g�*x��+oQVx�?o��Q�Ԇk)u[A���
�`9���vIVp7��
5 x�ǈ�j3��o��Ru�9���I�Rǎr�~�L��9#XO�G���u���׭vZ���|���Z�4r��!���z�ŏ�r71��%S�'��nҖ���8�aY�.4��m�׽>	���=9�Pi$G������4���M$]<~��N����b�+����c�`�r�T����w��OwU�V�<�F�b�*�����z�c����u�N���>wo�8��d�����[^:�I��:�V��6ZjJ�_0���F3	�*b?{���F���P��;��q�{z?e8���{H������,c��5h������f�;eVWx����<{�֭���8M������+��mmu|�@���o����I'���͞K�%���:>�_C��t�-���v�#/1����N���С�*i0��`A������Ĺ
��wv`}�b��un�j567]~&+�{�l�@t��]��np�A5��q��N��:����Y�ެ�M�KF#����rM�%bu(��\���<��E��(���?��eic�oGpJ����?Ó߶ݣ��^fe��k�Y�=Z�\��"�̕���9���<�ӑ��"԰�m��r%��u86i@��F��'�Ƃ5%l��e��H}�[|A��z�?���a������$$��B��Y<8��s�`W� �8����	ՋO���ʯ�l��IP��0l����x^}�5G1���c|,����2���쏎��6N ��6��p��'��)b-��\�(F_{J����E�����UP>��>H�����n�r���|��NU�HX�Wp������� ��G�HK���P�M 8~��1rƶ�{}�N���D��v�U���&��	��dU��0�ۛ5XZ�����e*�;|@��Z��%s��L�^ Y.;���G��� Y=%��{f�q�~�E�	�]v𾜕_W�D3d,sS*�qUj_�0?��RIAT2��u��h�� �X���Y��9yu������G�t?�ӖS@��f�������PE!����P�Z+�'?��t���A�<l��\�U g����w��u[oH�& �_�[�\�H����2�q���DǸ詶ɬ�O̰ΊY]%�c<�hӛ�A5`W���<�/ +�r�p��qe%Y$�֞�����~^1!Y�c��Sf�ԯ����X�=8�@�5���ħ�6�)� Zy�[�M��[%rX��<�8;;��❑�;.Q�m��yy��֋e��#\t(�6�e��?��+���0�����X��p���Y��*;��3��l�1k~��¬е>+L�2���ӯZ�L��¬�T�s�M31)(�/i|3M�q.$�~��c��g�:^vA��Hg	�w9
O�� �ʔ�W��F.J�BY J��-��.|c�OꟿX7t�6��L��z����)�~A����O���5f�G�5z��'�c)C�P�Q���cV��O�0a��F�!�a����q{Ч��TKz�K�~����F���M�jCY�#\e�1�D����P$xR�J<�)� �Y���΃<S��<ǟK�c��\���eWYz���T��ym�����r]�C�awѴ$��0�[h�g���-z;l#�h�X��9����{�ś�����c�����+Б�5�v�^{��A�A�ː_�m�Qѹ� N�}:i�����V��#ּ|��vrFXM��8���-�K�֬fb$��e���IR %���k����b
�����S_��O��L�VD^F�Z��J��ѣļo�*�)7���zD�v��m�S�|z��y���"�Y�Uj�6����YI{�T'e��}{>M~�W[�(�3��� ڥc���0 ���־����|W�rO�2��F1�V?6�&��֤+�eqP��3���Ū�F��ԗ�?�����Z��v˲��v��(����U��/!R
�J������,>+SB��O�?���Iw�U �{ݧ���M��W��,G��c�H�JV�k
�	s�>��'R��t�P���+�߮7�!����fZE)j����uEz�3�g��iT�ڔ\Qd�"3ME���l�%�!wS��J9�aEz�mS����V�Z?��C^�&2� �{�ug�t���M{R�
��O�	�8L��e�;�#����������_����tQ'�M��|wBO+P`�"kD�/9�Q��H*�q������ͰN��{*�P�:��O�HQXUۜ6
���Z\�?�Z���"�vq9E*ܪ�;}h���dV�k�|�ڊ1?\Zx8o���!/p�\n{;"�"�
}ڟ�P�I��Z��eX�Cuh��8g��f]�٨�򫟑����Q��yW5���Kuc&�(��4��q�@!d��|��V&C3W��݆n.�j� .�{
����O��]w�����{z�h�C��;��-<	W2����4{U�,ފd�v�O��阞� C
�l0u�*e
���u�P��qU�:Raa��jૢ�����d?��ԲU��j	�u�>`�e��VʞS7�D��������R��l_�_�r{�-S⡛N"�.�J�4����Aw����w����nxg����%������\����@���oT7Wn���p��̒Y��}f¹�rq����#L��}����:�,��-ќ��SP�@yü�=޾�#�}m,��#f9J��hi^wF'�Z+8`�.��������U��ݠ�'����c�� :$d���g���H�>+�(�4��nO2Y*�t�w�,I�Xp����[��|�ӿ��ͩ��G~8�O��[�ֳ��e�tQ5;7���/<�d�,��{��8	�z�Gi�I����Jh/7�Y�+��/����B�=��
s�|�Ǜ�I)��eFD��^eK����h����䞃5V,��^�:᛻��C$�`"��{�H"��f(��P�yn��	9֦�~��,C���܇��ӹ��Z�oC���_�)�LeX߮��4�@��)���_�)1�s��7]�{Ŏ4{�/�K���n���L�Xxm��~���6��M^�]��I-5`}1Ü/�?kq�@�-�4�ɮ�s�e�� �$�t��=`�������U�k{h��P7���)�9W��{�d �и��W�Q"��y�]�%�����t^�K�Б9p:��?%�wO3�Y��i���k�-I�\Σ=j{�]r#�ޏR�WF���2 ������SX&Kz�`�+y��� 3F"�#�%�s�E<ϓ:Ȯ��g�U�1��wG�dZ�TW����"��?|��r�kF�k�=v2����yƕ΍��@����ҥ�M���̈́0���J�����"��R� FM�_��Ĵ�ri5I���,�ɀU�1�Z��t�Nέ2f�e}h��O��5�����`�S�|�[�+c����;�}K�h��gy��"s����0*�+U��Fh��VK~j�xͺ�n�H'��#]����	0��/���wxV.������w����hO�0��?1f��d�	h�*i�+˸�4�a̽¨�|��KW�T�H(8 E�0X��U�e�i�ۤ+��¶N��>��4rg#���9=H/���=�x���G�����|Sl� ��9�*�'��K��"P����{E>���I-��<Zf��v��]?r�-�P�b�F��W�t�Y����\7��bm�m��8YQ�1�^�1�C�����[���D�Pwg�!��ui�G��ON�q��A����b? �l�bc�W����Z���R��a��^Y$�d���*����E%����^��}a%�X���V*uMz��{z����b���hD�������H���ڊ��z?�ף��a5WQ���n�UE�Λ>��C��~-BW���|u���vڛ��|��H�U���B欵R��9�wU���y���[��ɘ���$�s;�<�"Zk�H���-�GI-���w��m�W�~��}��ٶ�WBB�j��a�q{[�=�Bc-��?@/s��3�ӫV�3�d���|���䘲6�&s�e|�������N���7���O���J�n�gϏ�fx��ō[(��>|#���M�N8y�h�KXj���~�c�^�P�/Lj�i���~�[I�L�L.��yW�ϋੴ�d��ު�1HhQ��������>�46�"��Z��ŏ������R99����U�sX�|�j_X����]
I��k��+e��=�5M���t[@�A)+�ٌB������7V����hi	O�V� Ǿ�S�G�V`��pZ</��4�<��j
��-%Ye�dz����EW�ͫ�W�0�v��Q�L��ֆ���8JnX%Wd�X�7�6>LWL�5�=u���@R�u~�}�56f^��I=4��������W��������:�j�=K֯逍��٠De��5%
���&�-�v����7Dڥ���c��S�,=�z�EO�P��0.���S����*�������Cco5��^o���)���6�m>�7'oY�Ź<�����ZC�$)�k�}~�{J�xd��[�.MK���~a���.�6���U��;Y�[J<��<,TR��.�V�`_$�8.�j�w�rvg�{�+����*������}+~챣w�`��%�;�Ċ�cu�]���J
�8���R�P��������3Ge�Ȱ��@!Ry�� s��DK;r��������9�b��ss@"�S
K�BYe����S�ՙ'�xu?���
"[�}�m=h2ߥ93��� �����+���O�z닙�V�������j���Y��Y�=�_i�Π-J�{]��ңV5�m���-���~q,��7�:S�_YI�q�B�nzV�압<ZJq���;���Fo���4}$`;yx�>&*u���;Vޗ���$;jlo_�P1�v{��Y�&
z���qo����=[g.��.?�oĸS�,�|d=ݜ �Vm�Gkt���U�u�P�~�jwl�/��$�*�c����=��PD��Mr��c����AI����_]]$���&r��9�����]Bn��|	���5��?�����.!�^�H*H���w�*!:���akA��y��k�{���%�t��%.�UzR�4�qnC����(@�4e'�)q(R�@O��q�D��oN��)D��Lk��y�j��|��!����!��n�M��51���E�x�x�<ʉa�KN��[�䭩}��-L{��ȵ��&q�&/"Fv��Z�y��:-Q\]�īHӡ323��۫��H˜{s٦5���j�[K�������9E��ŕ����y+���C�PJ�[ْY���o�`�rv�X��(W� �yA	̼S�a7神ɛg�n(ty�Jr��W��	v�Z^%�G����'�����d}3�Mu��O��;2�e��4���.�;�>ƛ3.���g3E8T�.1�k��(���t�l�ݹ'�2�: C�E�z��?�&	�R�x���qM�nÊ,��\2-����^�g��!�3�w-0�|Er���A~�`H�>Y�)B�%y���]7�����IcB�8{�^|�S1@��	?����W���buYc��c<[8�¾wq������z}*텛~��[|Ӳ_r�Y4N@#[f{M�e2Y����ɢ��' c�(�?��%�b2��g��%�;�ݓ7xUR�<A���A%&��4�R��ȍ���kEq����3����Z���)z��z�3�*������?ASU�j�V�+�Q��(v$E�Q��|���uѦ!K�k��w���	�����W��-[�b����î���h:�@�vjhA�k �4"K�[�T9�%3p��޿�4V�j�Q��?�.�yͪy[0|1o]q;�do)۴���o&W����k3E��[>���`��3�͘���}oc�A�*<�\/ʱJ���I%t����F1t��6�q�ñq�[�8˨<���\Ə�0��E���5��I�tP[�`�_�M!�|�2Ukom���G�T���"U�Ow�lb����.D�X0�$�7�̙��-ewۅ���	��^.���_bd��db� �����������dG*��C�'��JT	}|�v����~	�g�P��zx�]5�r6I����:���;�W_�n;$� �i�3L�/����>��fQ��m���F��L������UM���)�z��s
�]��w?
�w��{���L�5S�b�:�>e�����Y7�/^������1m^�[�D@�E��c��vZC[���#ӫ�S7�#kت\���zP��I�/������ϣ�rr�סlq$KC��__�Z���h{��B(�i�W{b�}�;���5dg�Mg�?a��^�!��
��SM��TU�$t2�w˦&Ch����rL2*�)mNh�N\HQ,��g�Q�yn�!�C��r�xy5>�bg�w�Xi���<!��ԓ)��d�wSi-$_�"�D�%�ҳ��C��!�t��C�u0���i��#�G�T���%׵���X��Vv�8�HRS�Η�5�QL��X�[~�ZP�� �'�d���kKV��js���U-\�������@?Ɏ�=d�Rژ���^u�˯2	j�uK�7��������%���\��� ���r���\h�v�"�2{�w�Ps�0D\ ���{7�l�A ��f�������㪏�����m�i�]�C� �)/����).�׃x�UY�$~-�����fH�v���;�\��'��-�'��W<`Lt�r���tMz6��u���Wg��d�d�p���?�ѽJ��Z�{�wd_��a.rh�?/�[|]8�{�5+Ov��(	^޲���O/� �!����7
Ws]�b����g��3��-f�p��_S�)/�������x���Z��=�¥?v� \@�M�������s�CH��3!�>��%^��*��E��%�f�Z�٢�� Z�M�"=˭�U�q$��1>�O�i��M�}�Z�)�Uax��?S� ϕ;+�fd���a�KI�^<d5n�K��{����e��1E?84��[e08��� ״�I��-�p��o����`8u�?3y��@S0Zl�����@{
<����������_NH��/�lW<��B���vX�t��?�t���AK�C�w�����h��o҂�@��Оޑ��~�.z�!��6�5
�����a<A�G��B��:�6����T��i��t���]KD�>_�f��1|�s�������)�d��-����$�z�[~���<R$��ZH�n��s�a��\��; Ѕk��)���c�J�1���u�P����w���gO�Y�m�:'�����8��w����*�M�{�ڻ���D���n��iI����T�}q� Ӧ�2w�����o�-�Gf�=�g'e�(}�� �v�_��w����>7��^��Y�9�~� �%.����[>�����|�]�VGC�P��w��Q0|��X]�ol�_��|
����ߣë��d ��^��2�
�}��8�^��Fi�_׳qQ��_��� ���)ə[ټ��v��sgK��N�$x����opk���mP��Y�S6����܈���<
�8��;����.](03���S��.L��~TLL�Ȉ''g۴�^YtttnQ�U2#]1|����2�Xw�5����P-������={p��T��
��3�Qܴ����g��Re�{;FHK[�Q�i���oV0�~wwנ�&��F����׶������Joz�a���o�`�D���]L~�]��h�AO��ǔ�<��mmm�߾i@ e���Z&&��0�Ac�Ƌ7���qm��[�iz�'.�\�6�E��C΃@�����\*=e�&�����$�&&m+��FK,��b�:e�g�$97_�9�{��<۬ߠ��y����r���`�ԻFF��~5)U�����ԥb�_}7f���>����vd>�4�p]V�dڂ|x�R]�"����Vi�Rp�LVT�G���}� ����w���ƲՒr���u$���V�V����trP��@�v�M�g���[&e�{���Z�v�u�����r{�����>|�_J/sEJp��g����?X_��i6��\r	B�;��}# � ��Bש�U��������n|q��T��f��K'���5	�|BIk�q���"s�Y�O[DD��SCCce0/�o�_��mŤ�S��< O>v���'7:�����r0o�٧-ؗ��~r��%����r�ÅƏ��~�-�y�����Er6���6�8̵E����+|_P%1��~�,���(B�_^�<��4�	�g�E}��X^e H�����Sq�US'1�[]흝ZL�n9�[����סt����F~C���E������m�/C��̫B�MG��rF]��>vǌ�W�q`5��3kӯ�;. }���o�����xe��4i�jÉ��%�СR��!`����S(,rj��෫Vr��_�&A'�EDD��\���VT%��}P�io�k�ɻ�dd<\�S9����hw����Ax�uGs{L6�ؘ&+��VC�&zX��_kj��Ō��zKP�y��h-jQu�݌2������a�������\����@_#3������-u�^	���̿f��	��jlUUZ��}}�S�w��X��`�G"�l1<�&�v:�v�	|�yzz��pN����O�a�#ڸ%� �2�f�]�������*��9�@�{��w\�..�l�5A6i�T���V�r�^,�::%�@<���mm�ܜ�O�/^�N�/���c��Ȥ6�^ɨ���2�IĄ�}�#|�|�Lf�ok�j<д�Ti���yX�R]\����w��V6N".��T����V��i`�?}�-\���`��a�-+������f@,��Q�1�u�B���>���q�� 0����Y�Wb
�H����U���u�==�2�~�#����Nr�Sҡ\Ϻ/5 �3�_�2,s_7�&��}��󙙙{������V �%�7��NL��ϲ�I}胂�Yg/�����fŘ�W�M���ҋK|���SDK���BD�"p�}[�(�2 �+��J��� 	��-f+D�>$w�A�/�D��"�fBno���mmD#�S��ZEE�:j�m�"[o��i^�����bJ�R$�nm��CB�Y��:`��L��p��#,�
7D�������9r2�kэw;q��!�g�c$�k��o���O.FR��'�Nb���t>}�����[�?�.�wا,��R�������6�
��,�diO�HB$P��}�M`<�����`����(���YvrPDlJ��\��tVk#?d2a���k	�� �m�����|���􋈸�7�U�/��� y<'�]Ln���$ҧp,9����������:�%ݗDR�Y��������F�����{X	I��y�([Y�H��M�T�HH�.z���i��d���2;,.���!���«�+�.� ��rX&a8��	��V���Qx�����"��@�JFz=*G�p� ���S
o���z�T�!���r��[� ����{MdX�?$p�����Ā��u!0d�Z5�#OJ���_��F���3�
 �ZV��f�!���X���oS�ũc5Vj����u
��%����R�+'&^SM��sn (��w'�H�E�7x;��3��$�%KA�;:TFGG�={��m���Ê#-j�oɣ���7 ^�o�hj-GԌ�!��F�e���"��!�&�<�Å��j�S�n@���X[����x�1������0)-#���/� ��9ܙe��4�&�#��2�hg>�Xʑ���u�,�6�;�]�PUBW��v�G'�����rf,���<??�o������ɸ��lx�󴲋ֵ˿�Q<R�\��B ����Y#ﯞ��Ց����
�\]w<���'I(-�v!�H�!${o	7۵W
Eh�{s���q�B��6��{�����;O������^/�<�|>�����G/n��~��1*��ݹ�3�7[;���:&*ʒz��{�D:y�ڃt����`��m�J���i�yB�R_�R⮵'��u��+���ٳ���_R�btEW�(zs޽��)(�=�{�׫����K�Be�Qm<������b���u����å�x��y��֘�IUդa[�a^�f4��C��Q� ���; -�[�;�w���������~���Z�,����γYYYѷ�m�;D�k.|�����e������F�	9cD$K�� \�	u��;jnOcAd7����{�Y��8ǎ�޶eV�Q�Nы,6� ���,�Wo�� �J#�F%����
���ن�߂�DDd��$��z��ﾈT�H:i'x����*�_�9std���I�-V����پ��wg�A�c��wp}F|�
5a 	�ԯ��a2�w=��׎����'y�?Z ΃���.&-m@KTS��]YY�Go��XYB�$���[ a>�o"Uv��K���Cp[0ş�{h:���2���¾��Y�U�g]�8���rv]z��|��j�f�(�ip�#6e�7����?�w�I�.n4??mBQ����0m<"D�[�5;'�b�-贕匟���f&0(bc�:j	�r�ZE�GC��a�~��I�X�q;����/'@V�܍��Xg��g4w�k����s��пD�w�����7��b��F�����L�;���g���.�%qL[ޛ��5�+[;:�b���M���{U����@ͩ��3ri�=��x����Ia7��[n'�(�܈8�Z���С=��Xg%����-�)N5�	���ғ�I�A���h�5�򬑫Ą���!���299��r��u�9�����5[?�K����S����{Ub����J���"|~к�ޮ����Ż��:�*bG�b�j�8�S�+�l��0W�Vsf��!����p�!D���ȸ6..�ӹV0�F�����-V�����Z��LU�~�`���A6��#@��8�^]�(�� �'B�M����çކjn�!O�*� ��VxEM9��8^O�2�e�>�?"-�_���"{�(�P/X6����37F��E��F����z��O5p���ᷯ_u;�J@M�������,gm��+c�1�9p�(�π ��K{A���%��W@��j?Gsh�o�^�鼧��*[&�g�����E>I6����)����?r��oU�C�B	�W����۠���}IZZZ�Mv1]�i�"����~NNz�����7��x1��,i\���m�q��*������|),\�9e��B"빃���b�Û39�`\��p{Y���*&��/������;D�Х�р���T�R��ڔ9/��p�Z N� f^$����:at8o�f�6c�����
�U��l^�9�͵�䝣���K�(N�P��Bz��^�Ƶ@A������{Î�P5�wH(�}�^���[
:LI<L��y�$m�Lދ�֞��0�E ML��0�T�Ƴ"���K�:O�!�D5��][K����g��,Y.S�i7x���~9�g^��KI�wu���o'�n�<��*��t?_�ov*���m��<�8:���z:"��	Ɖ%e#5��df��r�r�0)��_�o7�F�ɫ�y������d���}B�7����ƭʥ����Yy�����rmmmXS(+��]B�qj��S��2e�i6��l�^|�h�LY�k���P�XK���������"�/H���c��e���f6P�oK���i�]Z(m.8���my�~��<M�߁�Y�3���H�X�<���H�R7u�Y9��&����u�0���a�)�z�Z555O*�2�5sV!�G�ymm
i$vN����m�~�.	���bICգ�#"f�c�Z#�vf�Km�FJ� ��sr4C899���M�hQSS{A�Rsk�:b�����pU���8��R��mس^���_�:��8�&,�Ui�=�h����$�)�O�c��,��ހ�6��[�0_�G8&�����3��d#�0�.��s� Mh7�|�T�����Eg������)qi���Q�;�ϩ�ɜ>��k���C>��V;��+�gc��j)��H���]6)>y�Y�m׹�1�����b��@���������.{c�b˒�"엽���5��ZA-����]�M"�Cݶ!�M�B��(�g��Fk`t������JW�k0����i�ώkڷq��;:I���+c-mZ���Lv#��`q�.�ţ[>T��I��4�{-��cM���Xm��x�}	�NL�u�vMF=]��ز��+1�n[5EF�!v��ߨ�[t�@@�LN�	)

�{-a����]I�gIk�*�4���#<o���a'��<C�*���zQP��Q�;���]=8�*/��/Y��IU���?�����n��s|4fp�)�ɨ{��6�}��}�v��;E�`%w��{���z���ջ�[Wv����+tTQ�����L6���)b�������_}ȿ�)͜��`k���!��/�dƏj�كD�zh�i�HNβ�sπ�na|oꓲ��\��Q���_m�2��>����>Ϳ���F�֯O{=����n���`�1��B(m�
����n���4ש����M9	�{v j���*Q��x�ć��I�?���ϑ�ӈ����ߏ�W���*^9�_.��Ȟ1��,�YN�ZS:}�D�on4���b���%W�珲����")�j+X��rMv�5?�F��K! ��Qر]_�2�Pb�(]|�h�|�]�-} �U�uu�k��
�~��"�K�,"@��Р�̆���.�R��+�Y@	fe��sY� �����ؾ̦QԘ���Ϊ,��%�?��@s�h�����+	�V`��ں��.�-��}��ƈc�<��8p�����U�����6�HUA"�k�ݎ޷����k���"��j4�\A��t�P պ]}�u䲔�»Β$f;��ӧO?��=�Dѝh[pڟK	����j�����aA�&��'��$��&8&h���ڙ�SM�'~�c`6e�B�cō��Y�����56��kj���.:戛��#l�5��Ւ�qs�)zU�wmǐ`���@+a�/=RR*�v^Ȍ�����du/���#�Ǵ곻�2�4V����GN�e�/����e"[{$;�s�:+��dpJգ�	��[%��3��K]����*����޶��v�&Z��Z��2���w�P�h\^Bt�3low�}�L,���FF6���)�߁�]IR��W#����P�����P�� uL4�[�TR�+q
�9}q��"�ed5�g�}&iV����u��}<P���p'��k�}��OF`;0la����3^U�����T���" �ԣ�,�A�Λ_��dk���f}��\��y+I�5#���N�oO��+m%	��4.�f�h�Ft~������0�XT�`8<��g�ưu���ݣ����:] ��I��tه2��Ȳo����
l%%�����W,-5u�:,��(�{'j���ס��/��
�[�^/��t~��>�ۣ�ܨ<�6�,�.��h}�a9�)j��ysv��Ƨ~��[BW5�H,�� |q��~S7�c��_t���g���L���ڌ��Kr��uG�{m`.n@����ޚ�g1�P;�n��*���=��B]TكnҪ���b6>�2H���dŞ�Xhp0�/'gKގ���x'߶�O�,fq���g�`o=C���>�͛�GG�ǻ�T{7a�F���UkE�g!,d�sD�q��U�r@G��(�{5����W�*͗�1[M�π��*s��n��D �Ѹ�[�/^ �ˠ&��LH�S����Ar�3 "z7;��s�`��0.�n^��j�q)��F�%Ѣ��Єn���|�m�4��ܚ�8�eR����)�|��Y����e�������K�a'T�Z���s=W��9�WY�hW&(|p$%�k_@M=��؇\P;���%b:iC/Q�������oǀyf@��j��x6M��Fh��z�E��M���ȗ����9m��oOQx��a���[���!��?мG&	��y�#FFF�$�,x���qD0�;W�����W��P�" �շuX�m��1Ȼ�n�M6��o`��G�J�*�_M��8�X��y ����5qw�n�R��T�,�F�=>�싳�X^���Au?--���l�?I��r��|��!�Ӑ|?�F�j����$�����c� ��B��e�ծҧ�(j�ҕݘ�D�H<x�L��5Tjz�ڰm�xؘ}�1c�ߩa���x���J�M�X�o�`�l�9;�ld��6;;{ 7.���9���;EV�G���g���U����Q�C2�붷����}���u�S���:�د�k��:&&I�a�g�h��v�7	TbAB��[w�%\9�~�6�+19s@��c������\�R܃��7(����CO��U�6��|O�&��x�y�E��~7[s���Z��Zh�٬�y_S.?)�	ygC��B5��I�(x�8�@E�C';��N1�B�l��»}�)`y�e��E���ӂ.˿����y�j��,��j��.���߽�c�T�R��v ���p����^��)�R�Y��g��{薅�R��H����OJ���%��[��)�wr��!�Y��K���];�����E�v_�QPd�����q 3�����߽;-GQ%�w���vs�^Q02>@;�o��>��}��8x8� �'�^|�R�Ԕ�/��ؼ�9�}�ڼԷ�V�s���y�B~L����g�c���ˬ��{�|]7P'�޴��]S��a�������#�_2��E�ء3��g�UL�ܳ�2�ئ!"��e5�4Q���D3�~�ʲN�x����:s�ZX��׹�ʛ��Z�.]�|��i�Cuz���y��

��%�W�|�!#�[ܷ��:�
�>�e����w�O��$$���;����JL�ׯ�D�^�M�qԁ�q8���{���n���^��tK+"a��z��Ǐ�Z�������w���W����ִ�tN�������c\�?��-U����3'`y��*ii��$/���F�0H�;ӳ���z�/�T�ljl�b��3��~�C�/wFh=2�"��M�̄so��V���b ��c��?����ה:�*MOO���Q���.K�'C��E�,y�ϥ����-XSG'3ݼ?א�o�w������cl���UD�,���[�[�|��Ҟ�x�{�t���0���2�}T�%M��������8�d�Q���E��,�땕iF�aM) �`۫�`�Qd��&�t�Vb�z����߳{������`���a����.ҽ�ԕԾ=ߐ��豌�L�I��)��}�?�N�	����t\-�@RZ�� A�P9Jw���ù�l�d��A�:������6D�2T�UTT�	xl.4���Ka΋C�9���;@b8t�ju�
DR��Q6q
���*�G��*g�l���:3�wi�F����\'�G�
-�(��->@�'8�p\<k'���,�O�5���:��v/���WC[���uYKKK`^��W�.0�E�mF2�o\�v-��w�ņ�!P�rܴ�8���F����Nx���UT[y+4���\����a�E�++=:ޜ��＠#|��SIl{�w�-A���|�zw���D�dX�f��yl��"��Ҳ���<<��g���	t\<��]�MAF:�u��E��P&�JÍ�i�����肂À.��EG�����M��D��t+	I	ᥪ��F\����[h+��aAA�m�-?E'�����@�qAQ�u�m�ݖė��|UlW��>��m�f��c5��%��)(2�����Z��p}��ӫ����MI��)���4�
\���]`����A�e%lߥ���[h<^h<�����l�/�rȵi^<3탆��%�Ut*2V���$q�L��w9Q�)��j��޶v�[���$����E�&׽�!�>�����w��"l$�MrJ
$y��δE�=Ӫ�Wd�.�/���:p�E-A�k77'7�B�1�Ǐ��J`SSf:u{�M�}GW��x�M���=�C�V��`�|^�~Y��$4>���$�c�#����҂���)��i�%~�׮��٣bґ��j�N��+'��Ԏ�-��N���w�b"u��rn9\�$�"�ʇ��|��lG�+��(ףlve�uƃ���\\���eC{�����s��GEd���;�ok��ԕ��!)4P�W��pZ��������X��X�Ѥ!c���bˡr����{��Sv��T�I�v��/�Ԏ�_��e%=|�p.3%t��{�G�lq�a�3��#��[f��}qڿ}ϑfRar�.�c
���g�O�YX؋+jjV�e[���� �gQD��X�Ћ�û��>��)�r�S?��jq�HW7+Ll�b����[z��Y�5��<.!���1���@�l�ޥ��gT�����J��@�f&1$�4l�F����sz��s�B�R�L�$)��"�8κԿ��4�깝���v��%=��6�=���	b���!��bl[��!�%��2L$�T۬c{��&���j�)�{*3��۬�>�;`r�(��Ήy�cK���+x����s���ů������vMM�VWW'�b�M^yi��Z�����4]]������WTB�(k��A�����
~�PS�������$ۣv�#�{�]�v��z|����|Ԉr����?&go6�gSXĻ��,�#��1	�C����1�Ko��=1���C�,�"�<��^���Q��6�{sa��VY�����-+�;�cJ%Ƣ]zMg��%2 i������������7o�:OcS>q:R�d�?��6ux?j�~��`��Xϵ,%(�aV�(a��u����Ei���S�FU�}��!_>|HZXx!�Y�kgn�4l������U��EG(�c#��9U�������$���Za��#`�P���*FF�+�M��&6z#������.�G���c�7�"e��*��T���D,�퇁�)�D��4�	������������wL�]��<�
��f�+ɜ&������	kN�Q2d��.\w������ ����������j��"��������OP��y����ln@����m*��X�#;�������n�q.׮+�fB�7++;�P��ر]����C������Rw��j�Z�s��_����$�J~sYVF|6�z��.���W�{�b?$��
�(|/���Sd��v ��|�)�{..�v�
�*��}#����[ۃ5�
	9ja|�����~=�7�؛�����)abٟ@V����/�y�n�
�OS�����&Q�i`vpp0~��}}n�eyLME%Ѷf����>����p�9Q�0v��ؗ�r���Z�Q�E��mB����Կ�U�Ri�F�;5����ǀ�z���� $v��8�"W4�e���!�V�U�uo�c�Сg \��y�i�\/�Wh���R$�?l��1 �O��MNM��pۣ�H@���	|C|��9۶?7���&-�7�`}
���X�-��;p����֡g�Z*�m�|V��iXG�=�0ԁ�Hr��pf����ݦ�h��7>��dS;�x$�&
 �~�o��ai���W����}=�&��\�S��! �2�sg>j(�����ӧ�|>�4�@�����YR���h��V���S~{�Z�I��]�\�y�=�̻sDG�8"H�N��w��|Z���}n���� �艬����F<U��ʷ�Po/Zĭ��t:;������Vo�;/\�%=�^'QR� ?Z��B��N0�̖�P��%9��r��~N�i�&�(%��N�2��9f�9V=Tjx�f��_���,yXaw��K���ٖK��S����7#�[�5u���ʏ�0�[=+l�RJ9-7�
�c��J�d'C�����-v���(^Y���PغǪ�F��𔑡!�����}��������W����R�K>ʕ�67J	5�^�bQ��v�U���Q�D��ꛟ��T�e&�HP����W��.6ݺ�A�S5�*���%o�����,�z_��������[�Rj��b��2T�V����������(SW��XӉ�`�t�ΩҁE�B��{E��d��x�C�������+țË<�'���X�bP�e�-��is�h�9:�,F������ŁZ�S&h;&R�9��/�}	5.�"�
Q���G�J�Zg7��Q�̧�5�A9e�w�f=)�5D4�1�Gw�/�Vo�e�5��ǟ�+P�31Pϵ���c]=�lB������Y
6�+��<D~���?��r��	�N]���rqeQ?����Fa���qW��hk&�P\(��i���VEK?��~�[#��]B��u�5��H��������	����k�����K��� �61Ȕ�R�,kNÀ��f�/%�Ӝ�3s���W&u~���u&H��\&tH�P��V��^[��g��Z7�s����P;8�]��u�J�� )��+�J��͈l���1h/h��|�+�P��7��67�C�6,E�D7#��Lo��ݱ�/���}/?�� D��cq�I�x�S'�\6���A�W�=b�L�L@b�u��5W�[�6"scՒ�?�c�@+�	0_&0������DR�fE�􅪄�K/y]��3.Vv�< ��ӳ����Lz�r2��g�Җ��Rhw{�v����"^� 0��8Ӧ���a2�Jd�9GC'v .�	���� �Ǥ�}��q��T��g�c~:��E�(hБG��Ѽ���"0>�<�j��_C'�7a�t�� +9��(J���<K��P��А�\u��g3jP+& �ul.�'v��VٮT�{4�����B^�w����q��#J�MO�eJ�yX �V��Yyr���q�/��F��؈�9�K�Ԭ�!���zU������e���WS�t��e��K��7�c<J��v�%E�n����̖�g3��<6��wl����($恼�ĳƞ���54>����� }W )��/:s_g�G٩(/��~&�K��`���,y\|�����z���94��7�qb�T����'G�2�?��A�lD8�E~;���"-|c��G����"���o`�o��셎�����Y[:��C�̫ۯ|��Bq]����^�2�>&ד���~�Ϯ�M6���lk��UI��_[��H�ыI�d%��+˞�z.���c>JE�K=G���������3���/WAÁ<gq�m{Y�QYgz%;�p�h1VI�R��o �*�%N=5y5����[f����>����=�&Vf`� d�~�����������lf���J�L�?�n�;2b <�9��;�7��L6�]��_���t�������]C�S��a� ,��cQ QXx�j�lQ�+�in~t�ܭp�թ��D�_�t���5Um�Q��9u��9�ae���óR�V�[f�tsl£�� ���:}f��E<�6b�G��]�(���1'���ݯ�� 3Ĺfm�����}-��Gi��%CT�6�_�Y�T	[9�&����I ?Y�Z�vQ߰tk�V2�&c>�)�����HߵW��2�[#�%ft���w ��q�9ܠ��(��(8�����V�EG��5�Qzzz�Z� �b6����`�{�����@v�_�Zs۱�>��k!��Z����K
��%M�o��>�黅R������!��a��.o���}4]\	|��@}r�.ko��0�i���{�+���iw�mta~�-�J�SS$_�8�!�D����`�	jT|�����i�-ɜ��4۞b$�u:xu%JX) �/ۓ�@�Cr����м?����B�
L׆�#a���6݊������!�8$�����oI�[�S�&��~���=�+l��˩i�f?�* �g�3���2���p��#K�v7�8T]aW�}��)l�T������v1	{���|qB���-_?2*3;�Vf���ğ��/�.k����>}[�@�)'���Z�x�EIΏ?v����)��']�A��� �+�*J,���D�B���j�j!�s�z����Dݞ���9�<�+�fZ�^�^�H�}��3;�a�x|�}fr�p��0\� {o���
����#�7G��z�}���9m��%4�Y}��4��b�5�����f�Bi�F�������cO#�뽻"��r� �t��DhY�*�,���p�V��H���|m	�j������P�i`�W�Go�:�,6]iF����`��å�m���zp���u��u�A%7��S�]P�W�(�%$r����m]:���V�r����zY��۴�*}��s)x֦���'b�Y��az�u$&z9���r?������G(8����7ZR�Y����Mmm ú����%BGe�<W���M�33�_��{.��`�7�=xB]��6t�[QG褳Q���
<4�7���_l���Զ��T�z^K#��&����y!l�<�gJ������18IWh�G�4��P���iu�C��9ם0򎂴Ϲ	��JB鎅2��<��r<���R�%=���2��*�	����j�Ӽ���N�;lMY�N�|*_�t�J���<�Va��
8�
m��yq�]#���>+"GUO����C����;χ�Y���h������p��<˭g�d���r��k��Rtw�}��ߩ�#�b��n�̶+>�X�ga�:pD��H֯p��������`�a�*a�:U��QNh�߬R[l�����E�M�@5�*�#������n�R�'SL����4�j<�e�����C�UC��ԩc�c������%�ѾSlGT�JCxf]Tzr_����Bi��;&~�{z��.~YC�\�qm��g1~�4k/cn�\�[�>`|
)�Q�s^��x}	�j��mm�DNNNUF& ��.%�X#�њffS'���+��E��w��@"�t�`�}��55� ���q��<t7�D��Ӌ>"�cbC=�0��Ah�f������;O�B�� }�Bq�~�(���%�-9%�j���(�E*���?^�,�%����$)�w�{�|���f�w��r��A�~r$��B�Ư:=˯��Cg�Ⱦ7��y	.��7�EǍ�	?a£X������G�UΑ4���]���(�����L�آg}�R������H��y���YD�OQ�=�JSdM�$��fq�R��X��t�'Ҏ�+��7E_��n�ݚ�����N�-x���-z\�>��l.am�*g�����Ȝ�Njj?~�m$}kl�1 z~__[C��%��@�V���k3�a�z��)�7��B|B YO�N+/�ٻ��;n�_����i�p�^���x�E�#��5+����_�j�;��ő����&�f�l#�wG+ѾЯ.{�ܮ�\���X�j�y&�|�~��[����as�����(6�������y�ހ�ӱ�'qy��y*~��f"�q;7�Wx)����Ů�P9�4�%>݉�Z�?����v���t��;|�+Y��Й�<6�&k(�r�eo�!,����Q�w�&�;��&�F�-�úZ�WK���|�2T�,Xt����4�����ҁ��dTn�S,���фʒ���ӕ��}n�H���Υ D��=���;�=m[1���]d?�3RR��pR����l7ujz;�1�	_�E���B������u�>]b���J&o�Ӗ�p�����4ߒ�!��?�N����i�U�?���,��
eK}�nP?�d^�x�Uh���G�,fS��������)� ղ�[Ĩ�:�ݒ�9�=v?n:�c�3��' }�jU��x� /p�P_�Z��ζ=1��|�W+h�oU� �Uı������e$�`����Sc����?��[iQ�]d%��=��^f=esc�N�$��S]u����.zV��9=�z�UU:��|��-N�~E�k����Qv?:�� l�\�L���hO�*��=}�KU��jp�i	%���cZ���m��F,��y����}�/����o�s�W>��U�D�gm�2�sk�K�0�Зq\2K�t̘�������ܱ�fs�[հ�֦���.�py��������'�����ji�� ��Ǆ�H�d�SWU�0�=���B䞄6Jn7~��Ҏ��k�4���3��X/�ϣetr�����^6�Eo;���6c���;Z^�.�7��q��0yH�s��g�������(�Փ�V�/��M����"������s��' �3���)a@'2��ݮ���)�Gz,��u�(���y����U�����h����ՉMc�|��Ryz����^�v�~�E:rc5Uf���2��3Z!�Bz��� �*ߦLxN�e�g����%�!�������Yo���&��:"�6`��Q� �r�Q/�*c5������Ъ��wHd�?��?HY�er`�	����-� �Ě=� �Z�x���@��xq�޺�(͈�%�g���l�j��]T�r� nc(L�?`��U����p=���w�d��c�{|��<QO_x�~�l��V�A
��;L��22������0���c�^9Q�mMҮK��~|��{� ��k|;���DS��MW|�!�d�%��?Y8��"j��m��xe�bǒ�N�vnX�Е,��f��H�'�-�ǜ��CFa��\���Vc.��1P���\�jB��V#�����?�b���h̦O��4��z	�'�v�ڏ�s��k�+y���I���&����J�<]$�N��-Ч7Z�ݑ��Z�^u�P�1J�MS�˫Hqux���:`d�=������'�]�m�l�w�j���$*���������Q��d|�G��m*������B����<��I�B����1q�]p�M8���IT0�h���i����J=7O�ŎY[!���@�m�����2c���s���(Q&*G�4ㄜ��yP��@=�+�/]^%�M;T[�fت_���8��-\��}�p�c$p�&�k�I��'��F=�-�����Wz���/�t�f�0���fѪ
��\����d%P�����Niג�s�{���Ht���{�6AwzB9Eb�NSP�!b�5�����_�4y�n��k ����0ܸ�(^ܺ�a"�,��0%1�&h�i$��߶G��gM���p��1��M�-c���*g9�^&�A\�����x��^.��|x�}���A~�R�e�}-��9����N��.��]�%<��0��j?ǟ9!f��?��6k-g�s�y�{�1�0�6�f'�V�Q�S�����1�,CY�C<�?���G��r��{�$�<>_m�-Q:@�y�UO��q�>�����n��ᠷn-N��[��)��,F�F��6G����q�����jLG�L�ۑ�q}���Y1��Gr�FT�
�����C���6wNۉ�L?�Ɖ��o'��y�������	�P� ClE��� %-��]������w,�;WY&l(�&+���n�v��L�F�A�vp�,���׭��S��&z�e�Ky8��,�fW�?R�!��>���Z��4��V 1�Q3���w�I���8��%)!�O�^8+�t�$EA�/n!kw�ū���s��0T�n>M2���O�]A��c D�Z����c�Ov���l�f�lv���j���5��4K�"��>��<]7�X`N��2���9�R�2Y����=Ҷ:dטa�-/r`�\z�>c<�G��	��ն��X��$/:���nf�H@�xy���ѳ�)*�
t�aF�<�;?�dc�����8�/M|:w��Kl���|f|��uu�B��W%��>�y(��`$�P�v{��ׄ��&)�孺ڀR?6� 
K���ce�ߑb�qZ�+�9GI��m/�팴BJVT'��
)����O�DK��ʱh_���'4#�tR���]IЋVO�='�UkG��k��4e�L\qV��CXﻇ�}�Ub
����S�v~f�Ѹ(�HP��>7�=��w�"���ԍj��HɖL2_N�^[��-�u޼�*;{�g��ͭ�G���F�+R��=jwU�t�o�3X����.��yUڠ×8�㔁��̮�sa-���&��Eb0O��}�>X>�J�tqo;���U�@�ѥf�WGs�2��%=�x"��\�)��/lӧ���-2��ur���~Lq�V�'f~�����H<�dK������Y5#}�mM�N�Bn����Q5t����y�5����2�:v2X�}�~�泯�q�h�n�u�e��	��=���V|��0����$y�u�-.�@���@n�P|�����ƼUҞ��GSXn��#F�ÚZ�*=�ظ��V���;��QB��w�-ߣ�b]�n|x��5���NG�{�Z㿧~���i�I�?߬2f�	���V��F2�dهu��֕�$����ˉ���/%�xR@^-�X��-3��SJ�;�ߏ�Q��٘�o$&;ޜ����^N��F������	��-)�;��[�;�@�G�g4N��� w�e�ŵ�ӾH���LȾ0[N~(�,JRq�����.��v/AMg��>,�N���F���\��C#�/�������2V^�f�����6u���-�ҹ>FT�NL�M=�!��������D��h�	p��V*|�E�e�b��#~���s����ĵo�]����r�l � �ɽXm��[@�]��E����i��Q�'g��U��.n���Cl>FB�)�~�����~�1�W���VK�椭C0ֹ{�㍇Rٙ��h�����7�F4M����,���yqJN�g�ՌX��/��8P'�RQ�nw9ŸV<���u��C|<	v[�9��?���y�u�eh�K�}wj&R��D���O��IRU���Ή�L;q�rm��W����<\�r��_�-����nr�_&os\�s'���F�]�]g;+}����}y�� �@6'��<�[�+T�%�y(�gI�p�_0���`�����b���C��+733>��Y��n��@$�M�����x�&�~��2�|tф�����Ƥ��h�r��>�����ϸ�fsB�P��8���j�	KS#��6"��J'�D�����nH�΋!Yf�i1��Y,Y�OԴ˞�v,0�����#V[�� 1�[�+�.
���X�'Ð�c�FW�$�⵳�}Pz���Ʀ���Kb*M���@�^t�uk�a8�=�W����=�T�T�D������>����?���,��v�@�`[GO��8�s(]�~��:r��U���v.~�θ�w}̘Ő���������A��bۤv\��ȶ����* m9��xOS��r}Q5!Hr)����� �n����^���a�=Ͳ��T��:�T�ǯa��!��3����n<s�9�;[���֝���ª,�{��K@���fɫ����C���_����?'i�g�b9Bڥg���m$�'��iM���Ν�����\���4�A��\ı���vM	�/���]C�l��'���&�_۰�= ��ZUs��hjC��:��~��/�Y�;=9ǜ�<$�r�����㬹ɫそ�f3/�%B��MN���E�D=llG���6w���.�o�m������,@xb�A`a缹@����![H��4�wG� !Ӄ��﬽4�w"0'����W�����j?�����Q�lD��������em{X���9t�-�x����A8v�ܾ�F���j�"�M�F�k^?�迷֡M��f���*X�Yi$ �/Y;j�!��rhgr�P�ؘ�x@;�t�����|�O�,�S�U��!G�,w�������Pg08��;���ou[`kn�c�=���&n�J~������.�A�.]��@YнZ�n%��坧��,N�Y�0�b(��g�=n��'�޻��<uG�Hn��醳]�kU�O&mB��Z������kyp���?���:,�N��N߂�t���DnC�Շ�����/�����o���~%t���GH�㷯�{���PI��ڰL|�$hz�L��9��cF�&�*'h��Ϛۍ5+��*�s��qf�2(J]�:�=ߺp�*�-2"�#���g|��P4���FM�&����:��=)a-�rsk)Hb�4�Lv��k!��M����Tç���$�6��z���׬��Uw2��
�ݟ�Cǵ��.f��Nh����g��-�۞��F�����Dt,��Z�x9�z�Ķ��-b�d��O�I��͎�q��K�q�.c��%uʇg��묬�@��@�w~cmM���}��!��Ys�s̲-��96=��[R��u����������N�2��!��ơ��1���(�J^?�@��\!t������[��%�gg?.���d~�r�x}x�-#5��ɯ����?Ӗ����S��Ț�Ũ�,�}w��v9�:MO]�+ҙ]I?�e����60��_�*߫�ʴ�<<��g,>/M�{�9\-Z����_�����9�qff�f�L�O�.S���0n8]|�	���Wk��H�{3J��Ob�o7o�����X!��0�O�Z�B���؉U(Qz����l���uD8Oy��T:/iU�ZC�>�6���G�m����[�J�	��t�E���4m��X�j����X�UG�e���G��\��~�u�2��)O1.a9v
ߣ�[w���	�f'����ure�z�ޟSu�N_h�L�q~����Y�L�X�8h��֋1��Q�!�:2��V_
-�'��I����=���S�啹���� .򼾩�2��5�ͭ�fx�vi'�<G����x��5U����J�$��>��m��&�����;m�y��D�4����;o ��}aZ�+��kɍC�onyyO'o� c_��V*"����c1�������4j"ﬦ�N�ֹŘ��G����
[�+~�3VWB��Պ�,��ȭ�qB%xR|�Q癙�s����weL��[�H������u������e�S�,L�hQS���|o�,��K�U���GD�� >���vO��Vm?Oq�!�,'bun�V32.�i��i�x�N:�j%��b���oߠ��%Fs)�S>�������-GC��y�4��4��x���YmP�h�r��U��D'z(�'��w����ln��E=ܳwe��jc��}gDW�� V!w�0<�I���ʟ�)�q��B�s3	���s(�1���7DbY����v^�b�H�����0u@��c.T:n}���W)��%UK}�S���;w�hK�c���rcJ�l��T'x����kj�����&�"�T�UQ�C@�H��{����;��I�� �H����z����������3����gf�=C4��y#ʶ:~��ŁXLF�&n��� �w��L���6﷯�j���Q���5"P������)|j�^`7�t���1Qu��4�?��ty��]M�%^���gӰuT���{��U�ՙ�s[G*M�W�dw��R�Ա�¦ݟ��^��0����=�&�Q
����K$��H��$�)d�u|8��nO�?'xVj3@[{@�^��(����</��/Э��s��h��㪮���9 I���j��Y�f�ZW\-3��vK�rgw���+peQ�je譊x�ʟ��2!͎}��I�}EB�R�ڻB� �մh/�2��s��.���9\>'����c��gmS���׏�o�d�2�f3"��gus���M�<��J�D�>�U��29�3���]�g�H2�怷N\��W�)���Ƥ��)sLL��H���Q^J+V͙q�&7�I����'!�I?~�@�qh�eTt4xY���U��+o�f�-��,J[ ʢ�8Dx_e���<q��<^2P�uz�{�t|�G��L�h����'�t�����*�Jݴy׮���/�U4��$ܬ�xE/�+�*�7�QU���N�XUOm1�9�r�S�Zmb�)�)��f`��J�:����Z8E�J����:�F�����˻�|ܒleej���`���ԝjd�BG�UO��C�������s8$%!��+����X�͢��0���2�sv�f
�,?%�FX�/��*��3�|�;99I�ۅF��*ӯs{[���Đ���}�\�>Ⱥ=4Ψ�����v��m:�A�)ѼA鳡J��\W�]Q��y,�Z�x�d������vU�?Vh�X ���`��O%⽸�%�|���]ɘ�t,􃲌� ��4�3�M8�+*�'��kq�oD�BO#+^�& 2��6�-f����6�.TbA6���5T��R�s�6��U����WR[���+�YoF��\l�sA�px�}�ϻ-y�h�;�E~�?4!������Z�G���?�x� =�cQ�BZ�aL��@\+��G�f��g�ݿr�?�o7Y:��)~e�������r?WX��E���1��X�����O�[W%̈́������zICcC����.G�[����71�C�^n���`CnV�k���O��f��ZB�������j���s����'������+�F�`��i���0��O���e0����LSm~cvK�d��Q�:6�_ƏqB��#Gz�Q�K�.vS�#+�O�������J�h'�K�3r0b�4�����,��a�:�Z"�r[��5h	'�wW�n�/�t�u<�o��1zU��㕴�yP����VZYA�cq�"��C3mpp��ĎǕ	��!E�I��d3�d>Ӳ	�p�'��!��+�L����Wʈ��O3�[|�����3�-�J���5Q<>	<���~K,ǩ�I����1�z�{��z���/��Tr���S��7��o�쭲-J^µh5��AW(�)A&�!��+D�A]J�
�u�M�V�ia�նuD��&���}I�Z�_���O�C`�B�=ĸ��.5�k�q}�;���
�r��ֆ��������]԰���aٖ~�A���Gܵ{���e9hW�|��ʬ�КtϘJ��	�wB��{�0\�+�rɟ��з7�')n���rݹ��{��Z�ں0^Ю��ݵ1u�Ý�zw���6P~�pg@���zyV��M~�}u
���c�)�S&ʣ޺aCm���n}[�r���}g{�_��jf�1�,�`ɡ�*!)2[��0���.�z�T޲����5���t!�I�i��V�e���o������{�]\}o��T���d����J���f�ӷnݪ�:\�E��Z��*Et>�/�Q�"n�v[hȟ�Q�c�L5��B�7a��>g.���'>4���''++��m�ݞK$X��]l��E�*�T'�Z_���i�9�j`��r���􇾙�mq��]�6W~ы2��[Q�q��6��������^�����!�С���힎J�k����)-ٖD���������f�=�/��.���eCf�wDz�1�A��$���5���Wx��du����\��K�OH�u���Ԋ����l5���Q������)����?ٿ;]�:@���ק��P7f�L,�b�	��o��`9����nos8͵6��.��������ҹʶ���A�&9�0�X�q6�x�>ۘ���<�E��$�hN�K����1䈜S����q��s��"��b�c=���%P~�0Y<��ݣ��
��X������lńl 	R����<Pgba���1X�N^k�� o^�ܳv/ehݘkX�
��h,빷���@���9�l0�C��H��Cb����;�q�eG�ݒz�ܺ��9J:���(	J)fx��,S0�;,��vW����D(-�z��g��_В�|���Mdr��~�fkؘt��ʫ�7痗_��=w�.�.y�P�-�V�,�J^K�|/x�Qu���R��.��9e���jT���?
\(+̩���5c*�߷�������>{�K��D����Ӱ'=�t���`�]#�����eX�2����[Ұ�<�r	�>���^`I�����sƗ�=f[�{�|�~^O1����N���:wL�j��vZ�7�3��><�g5�ZUSKCJ-�dW,Ss�i�CHѩV������ǁZ�k�O���lk��ໞ�ݍuNKJ�Sb���̨�Wp�9h����D�����/��w�i#aY7�.�m����q�30s��[{aS�
��6#��~�E���%���?���9P�@g��%�wjA�<ŧ��B���6���ۀ�S��Y�����sۘ���*��6�!ⱇ�!�;�j����D��R,b8C��d����K���k
w&}�4�H�'99���cr5���k�������B�������l>��Zs���	�V�3{�n���\���f�95��{��O��@�"��nq3=�gk�;bh��-�[�$�j��7o�^M�� ;ʼ���pq9-ZL�p9#<`Od��n�pֈ�N���@���y�����J�w����[&����n�<y�'�!2��$ep��0z�v����F>rh��7R�&�,��c��ce�A�`nM��6�nթ[Ӷ���ޛ�"�?h ���7^e����}����X��aVVV��o��3�r�L��=q����;�UV����~��+�����k�^w S�@�M�]oi�9��NP���Y*�A@�*Ѯ@d�����_c?6Wx��3�|:a�c�ѫ��~c���~h�[��ŏ3U (���Z�R2e�������߿`Kz^�Y�1�C�s��>�����]��0�W(I�j�/O��(�@�Bux;<5��x��t�(��~'K_
�=�/%��B��Ώ��G]������*��^J���
����.A�w9(�>�G�+�b��XX`�4lˉNݟ���axg���/J"m䇈��g��o���63��$q`�j;i�9��$0��fo������w6}��N�]��Ax�4v��؝���C�i�@4"0a����1�&�}��ĭ�����/���h�u=�m�S� �o�A��Q=��� �ض��G�sK���r�[��`��}8�}���\�9�Y��H�k�xM �y��8�C�p���kZ�������k��M����;����׻>���+&�V�q��U["�l��rj�,���X?h\*�eD?��[Pv�(]�C��[o�Çc)y�v{��w������d��U���j�f퍈C�L����m<���P��1�0��i
�r��'�j�o���u��`�a���������x�{��iNZ�o�����������oF�'� ���%�{�]����%�������PKL���&�k�=g���)�U��r F,�zUL���09ɞ����cx�w�0���V��������פ��i`ڬyሞ��ʉ��Ktt9O��	;]QX�E��+�9\f��[���:hdć�2��Iৎ��4:��7�e��v)f�G�gil�PUE��V9���͒O��������ퟟb�ľm�p�*�@&7zU��\m�꠫��rQU�#ߖ����ǅ��
F�I ҳ��J[ح�"�<y�y@�B z���bg������������朳~1�]�J�UM&1w��g�	.�WE�F����K�'�DSPP$Z����m�յ'Q�	�(_.��k�4�KdƗ&��'��r�~wd�S�Qh�a��HDbz��0��+���?7$R���=A[�8��_ߩE)�pF �R�P�lH��O��z�paxm��N-	�n,���>c�1@D�[�.G��ű�Nִ��:\4�-�ދ�l�OIztO2Q�������'��hhd�e)Y�[��H��ũ��� �^�B��i�!�>1��<AV9�-���(!�<��f:�>��}���;,>��O͠�F�"0ơ���-�q�#}����G�W��8�į#�Ư9�*n=�^ncOq�^�fu�@� �nPPeٱ��SQ��ڽ���uzH�A��(E �C2��*���&��r��y����B��z�q�O�%���_�mP����8�w�{[�Pح�v��.�	#�[�3�fk�mB�%\ۧQ�����A;1��
��%~,�� �C�t�D�Yw��̦���v��P�=��Cࡾx�� t��=	9/�����[�d�g@�3�G�֒�WI�-,����7�F�E+6��1��@sޝ�:+f6DG���$Yv�uV��c�ǀ*܄�j�mII�T|��MP���iI$�T�wU��:�ZP���\-R:��7\�_�Z\�3��2�O3%r�(	A�����b��P>�ih���+j�r�i�OQ��A����b�d��e��Ŧ���[�UQ���f��Z�n��2���Y�7u.�m$�Fn�D-�e���y�M�p4�����=��E�]e�jub-���`F�gGKK�2�QT�)D��QJr��#8�&��I?(� L]��s2p�9m��d���	�O�(��{��y������>@�e��;��� ��I[����UC�c��x��{k+��^�}����:�gAc�(����d��v�<a�+���s7Y��2��1�j��^�1��w{R���|!§��G�P	� @s?�q�Nިݢ&#3?���"X�����o}
��\����kjf&2T�Hkv�[cA M�P��[�v���E����(KMMjT1�i���b<�Pp0g	Xs��j�t��̃)�#�ƃ�߂P{B���Y|�%�H�Y�2;W� x�?���2+������ ��k�3{����βHL,-j�';���=A %���U�����s��Gj���{�'�����8׼@�����r����eɢj�oB{{XO�UY�Kۓc���y�b�b�^���q��w]{.�[+ϷXYYA#�a(�;f�'���C�p�,�K[���P9�,�w�2�{�2f 8|%/������}C׶���g;U��Һ3-�Due�iX�d��x��?Y4LU0ATl�W�C��N4[�]��vGd��yH ���r��@eO���]��
�օ�͛�&���|�{�D�����6nw���I�(s,���O���C��[U��E�2Y��:%FoD\זˉ s�	�O/�y^�ṷ$����J�j�c�*�Ep `Y�3� �Q��"�c���`o7�P�'$�V���2�] 'c?��GU{�O��į�ۋ���&�L�	UQ�J+
�r�@bEs[�C;����HN�9*��88U9���k�����Fl�o��@���8� W?ک��t0����{�xk�*���V/v̮XW��D�l��@���j�6F�^�/�է �m	�Oj��j���ſQ���X�2
i�L�ߠ�bg�����l��7m���h0����-֯?\�"�� �7�
�&��Nޅ��|��`�����o� ���rk"�y�����U�ꓶ��hoo?�O!'�߼�?���J����p��Bmߓ��;*�օ�!!�J�0�H����!�o�
���Ud5rlM���á=-�0}�%�Ԡ�(�ca��k�PD���wj{G�S�"�sb"t�777���y"ХQQ��c�X�V4���ϼ˻�$�&�p�k���s��J�W�s��>UI�������zõUT�א���Bߵ�6��ƫ�q�o�V��躗&����¤�%� _�lcz8s�ב{��ܳ���v�YA{}M������ͭ�܀���� NIIC ��'(�Z��Z�,���[F�gd�mEm'�r�*�È��8㦮�ۄ
;���++�c����ُ[e�<�nؓ/�.�4����j��wｄҷ�_}��/Y�f5���h��*	k���0\��p@��|��2-y�vWD	����%�_�4.��0z �E�ԡ0��k���jT���"q�[g� @3��:�ܢ>Њ���0�v�$x`m���,��8�A��`es���w,�b�����^�C,��C�9��~��8z��9|WѣU��-�����������bӁe>�zu�=�˔ǒ04o��+�_]�b�$�O�[~���2&!��lN�b���w#���qCh��4A_��>"��,�R�/��V�U[S6�̽�ਔ��p� ���[LMM� ����uA�-	�E� ���T�(��?}J��������s�V��-v^^^�֮��M䒝��Eae��&�?���!k�o�#���9�p�Z�S����J ����:�V�Cg�l�w��I����j�N����G ��Ĥ�����\� ~�OY���,t	]-��,r�qT�^��K:�R�vq��	��v�A�+B*�����<���sY�u2O��<s�|S��jQ�1TcS4r���N/����:�5�9!}�����P���ol�c|pJ2�/����u�ד���OJ��|�����w>eC.P�ڌZx�f���A}ay�= ��:/{��U]�"u}DD�����>�����{���W�5 ��*�Ê�ƶP4)�S�p��6r������עLP����U�j$S�T�����i�?.7�Ѽ�N��n�����0�[���n�?�:��9'��h_�f&�����U��X�b$&@�\�!M__� |�ٓ��""B(2���5+���t���h�Z�1iU|�lY���z ��qi�TZ.T�����4=b}��`{Q�_�z����]���F�eD����|�x���3U1H^nav��PUn���d�����_j"�T�|p{�� u�F�$'3�v ����ch��Z>^�Z���a�5��y֩s�i=�
��o��P��z�W��]�v$|�(7�c��ƨ�����W�>�������l�v+�F1�[?Yk�w=i�8E���B!�֢5Qg����_��n���U�<}�
�T����'CW��X�z)ovi�Z�A �JO=�l8�͞W�S�<5�V�z���%X�w*���q���Wq��p�.�WZUN!̺�ٿ�J� L9g�V����(��ѷz�-[�]��A9l&j�j�/^��;�8��Ƈ�s����ez��A�f�䛹���P����pgm���^ ��F<��1�q�C�����	 0�>��$�B^�q?��M-�B�r���|��t�=^���%z���{�5پ�Ղ]�ĄX����1I׵�T��D$(IC�7�}�T1��2!t�� �v��s� ��u�!L����o-�F������= >�����p�^��W&����}a��_������Ar���9���N��<�@��lϑ��(��q��?��cx0B\zė�N�0�<�ˁhM!�NH���d�a�2�	�|��V~a��2o�P�y�G=V���_���RH+R�9�����m��?��=1����Ejs-�x�}��sz'j�|�L�(�v���~�����R5Q�/��s9���AR�W�7�窆6�ȣ��֯1e������<~׶i��������`Y�0�Y2��( R��yO�{�X��f��"!=�G 4����CZ�E�����8�V� �0���6t V�H�Ck|#�_�%�_I��fgg9��y��M­��(bo�
_A'�jfΤ����Y�S���Ҷ�Qof�^��wQ����=�"w��l�འ��.�Uq�<�"�G�~��5��2㋑b�O���H�����Jp���q����.�&&̩���PT��Ph~=� h�,=��/`5*DL�<��N]@ɣr����j�3Nd�#�����=�6�֫֣�����)��Ɣ�T�ո�J��ك��~�#��Y'��]>��:Zj�$�m�|���*��ߟwA���!��:v�SK�ڜm�_$��ځ0��t�PFn�O;Cӥ�%����7֓���$�E�d䢭N�TJ�7vG�V�x�Y�LCJ� 5s4��+�%q��m$�6��	��E��{�^�a�ӥD�0 ��g��E\]N�GU��0�w���E	=�U.�BMMͬ=��V��O�O��O�18q�����:4�n���|g-v�O��C�_��������2�M[�j����+>��2� ��5`��|f�*�D�ӻ�q��0����>�x�$�����Xܣ�bOv�v�px?����rw�F���O���_q���;}�֍��@}�WP�Ϡ�u��VпE$M�i+�H�~�| {Ffr�U��wrI<m�ŋ�I���F
�x�2�٢ퟚ�d�55B������i���7�F�9�`�CϒD\���&�h������$n4��߶�� �В���/����
vV��y��瞓�T+�i����������vK >��	4/��������|=�ң�5�
F��O�����.u	�U>��+�^V8u�֭f�	��e�B���*z�{$��O�0UH�֖��B���-i*[1ADY:wy{PO�\�۝'d�c�ʥ�����[��%�|@�Օ/T�hYp3�E�2��!�um�A�q��D�����p&X�[������7��f����3�X������%�"F�H���=e�����r�y7cW��:@�SRa�\�O�>�V N��cgjb"UR���Z���uG�R�\� �t�n �bO�:[�u��. �31���-\����|��������>	'q�+-W�
�`{���W����c��⫅����XΜ�n�� O�/�)�O��r�$Q/ʨ	����6T��w��	V(H���2�Y85�s/��Iɬ��Fppl3�b�ɨJ���r�7s�s	��f3�q����;����B����l����S$6%#�}��T�4�;A,TT����"]�v
i���.V����r��ol���������())�J���p� �_�7�t;�Bs���i�p˕fB����uxn�>����SZ���$�ߐ�n����s�i�51#���ഭ��DM����)2v�i�eD�f{�K��s2��l���x���a�X|��/�ͺ��M���{�#ۑtYʥ�����&Q�e07mBP�չ�z��Ý�|
��4��^��^{��w���鵳x����l/DtD�I��n^�%�V.˘�:��{�����u�F ����>-a��<{�������y�GK�ı���w��W��F���>ay�l�����B�|ij�����W���A/�ʭ`�F�I��$�_��Ex�����$��B1f�&m���H�Z��m��e���(%%jj�m~3�}�5]l{�z���ǟ܊o������j�z}��A?�O`j[��f�[��`�?>A>���A~.�rh&��f4o�S��SS�K,����|�yxxP�8"��DA�AQK�R�Q`i� e�V9}�4t����S���=������,m�b����"�-}1�44C^���z����� %�k��C��{ ��(�"���u�^����|��
������ߺVS6�Ľ�L���,��H�C�(��k��5�#ҫ���=	�=�}�(��;{k��m~@8���ӧO��ʶ����m#n��:5����)y��V�k���vצi�#��`���,C?f�"�s³'���8j e=�A��U�A���\��t�mʣ5o�.���;��>u|Z�����yb
tp�^�`�r���'w'�6�gɝ�O~�����Rwҟ"���E��j�U��+�]mΣy�%(��d�8<Q`Aٙ?�yS��GOվ�
�S�6��Ҹ���3ͭ[��.6^a�^������2V/����Cou�#�@�U4���� �HGN��wƦ��Ez�q��'tH/���PR���/z�ލT�e�Y��4���޵��şw�|�U\�T��15�w�	ϳ��,K����'�o/~�,)�7�_�[l	<�$9-���v���w�.���6��k��0�<�"��G��T��% �⳧��ALűsk�{F�INr�=xQe O�=�����6���4V2�q<_+�8���4꓌*q~��+�S�!��>����p���k��S a���g�4����S�y��AΚ �ʃۜ���6��.�%��$hĨo�8��y���[e�q�$��R94i��e�_ש7#E�9��
��K��#�Nl�Zj��I���-7o���Nw ��/
�j9+��Q'�2�`��ݒ��Q����\�7W�wm����>�4����|����JV١|Zd5(�D�V�_�����$�F�]Z�ׂn��4�Z���־5�{m���T<!���0�zg��C_Aߣ�Vz�?����`�����H	�6Æ�enI����0u��y��_��G�����o��������V�j��b!�.�?$�e1Є	P��nӸ��B��ؙb/�)����R���G9���u)� +C�a��dy��S��m_&ݿ 4D;�J_���~�[��٥�j�S�qFUw���u>�߶�R�h�K�n��ñdvd_�U/b�aqI�Q[}���AH���B�^@F��*l�V�E�z˄�@��n+FyM@9�\/"�cQ���	�RArՍP4���M.�c���sr�!���XAY�Բ�s�~}����]0y�Y!YY|�ϰ0Z�@��� 5#�� �d�W��#���m?��}S��({R	���YÚ��|��:�:��~�"����f�Ӗ��.�A����)p)���onv�>�W7U�N�x���Fv%g�����Rp����Q	m��0U�,��몾���e ��L�����h�h��X.�n��;1��5�C�(竳z��'�zG���
�c�N���wd��F]B.����y࠼��6�Ϛ�H��~���\��U��kpm`*.��6α7�ƦĴ7�%܈c����ͳ�,�|]��X�zx,��Q�e��]"�/k��n�P4[k�-wq-p
��u��B��B�wP}��sr+�&��U�YF��Q��2�Y���"=L��A6�Q��Pga���*�e����ЎK�VoL�ho��h�>��x+X�&�܃:�B���L��{77�z��h,�oۭ���*�H��luX`Q�^ˉ��zZO¹.��uӗk�C�p�	�Dq��;nLګ��졘�+���^�
V}��5�<��A�#|��m���'8W��>ٱ]\7��}{8����j��B>�^)����\F���0���Q�K-��}���r9��Z�.�6QN��Ô��*�_��(�k��ԏ��͝����VE����ſ�@��W�Tis	����{~Wű���w��~D[i�F�L�z��]��{�ua��p���W���8��U?�;0�-tOe��$k5UoL���t�I;I�5��}�j �r�sn.:T(k���2E� p�Ptt})���<	�a��r�#����<ff��I�fi��*;���f$����iէ�F��C4��z���څ�g�UC�q�!����Ҙ�0� �)�5 �V��D=��O$�tK�/#�@-��oy`�y��)7����|x��yc�JS59b�1=�%$J�P�CM�yt��h�4t�6�K�X|�n��.x�Q^ۊ�Ǵ9%k��)���U�P��IM��e��r���5���g��'Ǉo=+>��y�=Q$���t��/���JUѾ)_�~׃�*9߻��Zk�Q���GDX���x~����~����� ��j���Ifņv����D�ԨY�jX0��v�c�W�%�
=~��y9O��ʔ�`�u������F�6�D~�O���ӕ&�$$�g����Z#K�eȠG��ˈ�Av1�~�G"���j�a��LN�Z�y�X��%�YOL�oN��kZ|�0� �2��g����c0 ���^fJ���^{ P�G�m�œ��sS
���~�[���ғ3� ��_�����i?��S�Y��6H8;/�;Գ畓?{m�-�8�y<� ��_�е�?����$<54-J�o��I�7���7{�&A�0rlv�侧���Z�5���50� hq#��&\��e�O������TF�׷�wr��� ���^)Ȼ�g�v�OW+to�~A�	��ٝ���-6��2`�d���,����K�@4|��>)���˹�y�<�����/߿�~����>"�V�^~;�o]��F�RP��X�:�|�^S����`���X�
r��+[�4�8U�M5ըN������S�96�d��G���rW�0�&���m�I���^��c� ��T����z��+������D,*p���
�%/Dm��K,�F�F>��r��$��R�M�:�ї��0��S z��K�~ 0�d=OAH�E Ɋ��������޳d6�ѥG�#���b��c���|3���0]�q\Z�=o���PS�����V���qKn���c�x^��M���t�����������������H��q���kN��or��v�9a�-��F���1W��Ħa����D(RLT�`��ߧ����z/�^��&�'D�]"����V~��� �z�DV3��-����|w�_ƃ��\��oP�g� d�
*��f�,(|$e�hT%���5����q����.�MFd*�|�"��Trl�qZ�A��pH�[;~��͜K]l�פ6tѝ?Wq�V��\2^��N��\��3��XCMU�X��i͸�:N4=u�N�Lq&����`ir�$�3B��aq�5��ѷUN����;�w�ì�?���E.��ܼƨ��v�/�?%?>���I�!�4����#f���Q�8,V'������k�=�؁����df	��{��Q���]�&����]v�3����v��� h�Ɲ�S�����.��	���q�:Jg���t�lҶzAE��PC�QY�+/��Gp��� �/�����u\�g+2}��j����ΛA~�^)UUUyy�H$F���.Ƽ����r��[�����Z���!n�p޾}���*�bڅI����q�O�DA��K�u~�=��y��^H���:b�1j�(!�˗�JedX�/qB/�I�ܸ�~!�{�-6Ũ!�!��a��z�1T��|U���F�;��{eI�����bm.YEEg�e<^	��:�0����|8�0Ֆ��^'d�+H���!�&Dj�F�t��Y��Nt��nY��'Z�(颿Ʒ����ڣ;�q/ù���[>2����~%O;	�֖gnҊgD��l1=��Bxi�uC���6�#��KR��uu��"�[�k��ٿ�fT�bx jQ"�g���\�J<��sIS���.Ӛ�@HJ�Ed�ó���i_xY[����H_yaa�Ѹ8X;Ʒ=�R�b|�;�;�>��L��{��'��e���f��[1���b8�]���lP�eek?�- �&�}s����/�y9�ک�p���{2��p�����h�)����9; <l�.)Q��s5��#�ӵ�R����:$��G/�O=��)�\{)��� ���:%D���E\�Zg����a�P�2���q7{^_+�z=��.�g���f,F�����*v��UX�@^ �-�rܯ�6�~����O��q���n��;x����	Xu��SkG�,`�E���Œ�T��C�e���T�;Z���/ڍ�lT1�O��A
��b�OWP���/%Dj�e��ZD(���H�A�?K�ҝ����:kDrUt�6,�	���h�ؘ�EGn�;��l�\?S<�������W�o{���`����&H�y��R���mel#�Յ3߿o���x���S!�2~��(���}!i��aÍI&�ó5�.eX��T����3�	�VG����B��c�g'��>&�bVONa'�]��"��L�0�X�A3	�DE����Oz�9�9AS~����'������Xx��~�Q���Q�]���1�1������{�ʕ��c>�P�|��/A�>�C�*��/�Dmm��+�X�[Ƙ"/�t�lo	�OPTx������$%��YI��Q�5�	:4��i,u.�=�,����<J01l�[F0c�1Rsj=��%��&0��F/"���x<����ٔ9Ā]}���?�Q��n�Z�MZi��q�bB��7�	I��>���sz��oќ���aJC�������"T�
��|.�����ΰxd�}1��	�A��&�	�(뮬�P��|U�5��E�V{���=��zZ�� q�?A�M[V�O��B	�E��7W�����
V�WrE%2��D��cU����w_#1���b�5�E��K�6�%
i���t1H:r�c+�ԕ��*���(��:�?��h2}_(POm@�mn-�,��p�G]���������+�V���H���=$���Hyd���.��ޠ�!
J�>������Ò>��VU��ѯ_�e�k9�!��)M��d�=�il�c	c����HYf|�`�kg��|3��2�#Vƶ�z�ᤈS%:c��Z�8L����L����}��o�KI9N=B2�דXL�kj�q�>na��L������;�J<��v-�W��S�T�v�iӵ4b�;�^���{mٯ>�Y���~��/���{N� �J�+0m?��m��߉��k�KY��>���L� ���|�aG3�X��g�tfq��;�A�Ǡf�@;Q�̡��,����|������o�a��%�mX�vةVz��t �2[�VY��F���q�f[w��0��G���4T��p�dӓ��<*Y�s�7�]u����Y�5�-��'<�"X�-v�G��Ȗ��V
1����9����\t'����Փ�fŕ||)Z�uϼYC�<>N�]�߽]����cz�s�N��{/Z���h�}�Bh�<w�2��Oi�U&"�W�/��mޘ/G��D�
I*�_����U�4����o��FE��W��]���eNTj��,�a�v�H8}�
 ���C���!s+��Ay�G�툟�򛛿�������|��Ke��x�'��٬%	)���gᑴR�����Z�X˩:���:���i{�z�w{_��w~.YAc0��D8�Bك\V}�ܤ���_:(��H׷�J�0D�����N���:��փ���k�Arx�Q|{���� `��[(I����G>���if��+�l���Ͼ��SW�1�?m�s���7Y���%$O��trHLx��v�0�c�`0E��i�5,1JX'γO
�%��>��ǃЂ�`u�خ��B�wwF�;����xx��P��@���W�HGE�y묬�����h:�3�+����X��.�) 6_��-��@r�=$$����"�$4-��`ې�Dz���Z'�Q�+tcg#��soGB>4�ܲ��}yš����������Ky�,K�Q0�<�H&1:�s�'�Ozd#�Ʃ�`�����ZC�gC���}X��97�t��n�4N#�m�ҝ���8SI�
�`^8�E�`��)�*ib��H������Nr�O�΢[�n[�~�>��Ky����\<��@3��o�5�P��o�E����yh6��7Y�.-4ހ��j���a�һ���$�1���+�Y���;č����#��1�����q,l���\�8��yR�@��NR@٣�4�T���Ff�VYGdl,�#w?�M�1467��'o(M����K��P�<��";�b�47�H��i�s§Twy�[���<e8-U�Gb$�R��H(�nDfDLX�����IsKȬM&ެ_E�`T4��]��R�н����&�ݾ���Q�V��;-����3�Nx_$����e7�X�	gzP<0�pQR�ƌ�~s��H�ĂO���	/T�.W�>���@��3�(c+~�P�=���������"�\�o\w�	~�־�q����M%��Ȳ�����Nv�f9..��11-�Q#lr��*���	�ADAޕ��ϕ����s����:̻����ݼ�d=��d��y���8c(��7?Gɥ��f��)^�,��ۯ�������	��;S�*a��~����:�q�cU�}�T#�ԋaw����`�W*����^��7	�5tWi�Sl,,B��O:q;F��}g��D[�'�y~����	��&�uUB�a>����	#tE�y7�	���.��ؚt����ȆR1,{��ea��1!L��T��X�������:��"L�	zP�/�?!�^�~�+u��}���;�]�y�)S���v%}�;�lɞ.2S8����M�;L�Fp�9c5��գJ^|1�������R�G���Ȅ@�Dy�ڶڑq���+I鶒�i�������l۟+�׻'��eT�*E�į���g6�oDw>J�92J�$�n�$kF��.�t}|�[�N�+Z�R#�x�+������0s�f-;?w'L6fi�������"�E�~��z)�3^+�J�����"nB辛����}w-����:Ϋ�����C���PW�Zφ�=�^���d9k���3o��y&�tn��;�����[d����T�0;J�����f�a,|�������!�D�j싟���ˏ$��f�-���D���dxz�Wۏv;�I��¦�������!�o����~����LF��^�t����:Qfߌ*<X��Έ�ߪ�(�Ҵ����R�;��
�
L�y�/�LF`�_��
�U�����5{7!$���D�'�ͷ)c��.���M�����s,���oO�D��q��&}�zBi�h���!�����%;o��<?{B�/�4���P^xL�����*=5�D�B�U�����L�\�ux��r�����߶������I]��J���E�:��(B�^�ҡ�|a��y����[��w?�c#F��Y�mG	6P�zW7�$��O�1�~"�*|?|ϐ1�&�d��=O*1q���G����wp��sg<��zgz���c���ܺ��I�DA��� �EO��h-��^��-zt�c0�F��D�uF'z�Q��v��s�����{�}���kݻ$0���Z��}��U�0;y�?�iX�k'S�p:�����`n��1a�b���Mt!��qحv����;.��7��j?�򵨯{P�pI�<<��$fWq��R���ROA?�.�QD!�A��~���*1[7*��\��3=�����_5�h@ ��ϯ�dӋ7?��jbZ�/v<;>��۝�D�gc��D�c��Z�#���m�IW.���3<�,��>2����{[�J�i`�Tw�2��0|Ϭ܍�+!��OO*X� �=[���@V���t�y5����eQ�|	'�,yǖ���:�&���T�y\�3S�3�n�ఊ����n2x~���:%%��,��w^��Ą(ҹ�w��O���g��}���H�Cز�]B���b�ÄM*�V�w����}?��:�Ew���D@���� W,1��H��u�:�q�(~&1���]ۦ~���+;���B��Mߦ�/����]�w6�ڏ�-���� g��9���*�N]��6yb�~# ��������Z�S��ut�=r�`	�����(O��5^F'Z�S���l2z�v&t�|$�z�ڐ���Ѧ9.�c�����]s�/��ʴ[|��vg�5���T`R���9;ЛEo�&a�G]�����$K�QUYA����k�U)"�9�]��1���7kF7c�����7�"�W���U�b6�x$`���-��g�$h�S�A�J���=2k�[�h�4cm�������jK�8V��Ԑ 
�N��`��K 	�rl\I_UՕ�8i�1g�FI�VeѿN[�Y��N�e�J.˨r8���XtY�-{�5T�uko=��E���0��kU�K�@�v�'g����f�$��]a4g��&Ȕz�"J�%��.�f�j��>�~�I���F�,��+�D>\��QӤ���*m=�<8 D��D&[A{������{�e����O���#"�v���t�n:H�Q���9P)���#Oc�����*�90;u��|��l�wm����h�eҗ϶�����ӊ��7Y�;䉟wG��敮U�{z2��@uj�b�3�&Vx[n�����p�{w$O/j��������6��tex=�L����79����)�=T�op�
��|���4�d4K��qf�[%N��R҉¬��um
35���_�y�5�|��ɫ�>�U�� �����ɖ"<E�v��V�{a���۩���;U������8�h����H�MT�ַpu4�sHc�|��L��=��JCK����X�ٱ��r��]
c$�M~�Ā6�!6�
��
ă�%/�T��L[5���\�Ƃ���o����"f����fWt��)#��l��9 Q�l�9ܛ�~U}�r�Ԅ���}�?'���X$5���SEU;&�3ؗHy���r���]Q7w�!��������+c<n�u��w]�r1ej$az[�S�@O�:�y���RD�e"u�6X�:�	�1���ސXN��Z>-�#�~�݀�i�z}���Xn�f͒���_�V���/��P^y��K ����f��L�nfZ+o��i�b��(�ۃtU���E\b��r7��JŢ7��wÎ9Sh��,5�S�R ��6�Y��"YM�z�%NO�N
��A��HDS��u������s�h;��to�VX�7�fg��(I�g��R;�)�ih��4��*>��+'F���̫�~%��Z����C3˞�H�����ɫ#��g�#7�1��3��ͼVk�筽�Wk��n��*�+QsdJ�p(}�m T�}0��K�:q���n1��Z��ݙ
�U�$�@����a������3Q�HD���߻Z���f������W�0�iwf�.�n�j��r��!%��*Ҷ��_�>W�y�ك9v-Zg1���(��k�㘘���z����o��2���ribf�o`@�-#�g8PQr)�m�s	J�F��h��yC��4k�g�.�1�:/_}`�$��}X�HF�͏��'�󍭡Z����X^�YJ�,�2%OG�H�(���{<%��r�u����04��/{����~d��#ãw���u b����Pf}P�F��m���Ƥ��}��Tj���]�]����d�����k�V����߄���t;O�ZI{S�J/-ӂ�$;�~�>��N|Su�,%�8^նe4�Zc���Op��i��|��y���4���o�S��Q�LzN�3��x�g-��c�<z���*�'@���;O�����c�o�})�|�v�ÿg�Q�ou�8���G�=&��k��#�1�]���I��ᖩ��t\�CK�2(˫C��yLs9�D}��#}�E�gx����;p�a` ������7���=�@����4JZ�z�r.c�n�R~͝\�am*;-	����q�x�a��ħ%�3}���ъ �+me��:ǽ05KV���Z��o�f}�ם"�~�u�`ޓ�����T�j2�X���d,�>J�g��b�O�ڛ�2���١�bY�h����ʇ<9u�r��p6��5�A��KwĻW�jXÒ*�u�P�+�,�#�l�އD����NZ5�Ӏ�L�J#�j�(�EuE�,@H/�FM���ֲ�uow���p�F�!����h��}^�dW�Uk��X�Am��Wo�gnY�/'N����6{�����[r�6X<h:�4%�-xm,MX��Q��{A�ó�Io��0aA�����X�e��$�{VyUNf?�M[�!���C[`���!:7]�SF6��,Z�_�'E������Th�6z�l�Ce֠� ��Ǧ�2��#>��3Y$��.f=�)"t�l��Z#��e���_�c��g�2i�L�F�сqt�İ���9O���di!;���t[4������qkwJ�F��` ����'��N�)��Pʪ����b`��|:!���Bאf�t="6Z��m�8%t^x#,#,(!!�:<������5h����8Ӕ���,䂹Nv�v�*=�4����Ro�/J���SEg����o�pTEYȇ���+�'�_��)��t���;�d�
R��o��r缚*�R.h7��:��mQ��B�USo{ېS��aaG`<����p�r�6��rcy����m*)�3�x{����7s���&&�tc'Q�����r'�� =����6J�ז��^��!~'9j+���2����8�ki�w�ao�j6x-���J�}c�.���F���Y�E����3�D�2M�0�s�V�z>����u�����v:�＞�n[���i��ƨ�7��ۊ+$���1��ER����P�:�X�J!!��-��zy��T:NT�ah4zo4I^�����v$A�.���x,�z�T��P���*U���p��`���Xo�Açw����We�M��ѻ vY��ߒ��]=E���bo���0�ڨ'6������fI��$ċ�x�M � ��~X�jI�嬹u��yrg�v!h���nZ�OI�2�z�g���{~�B��r��O�t��])�:�۱*�v$���cNY_�����'?�\M�;��.��V��g���@Č�<6�7\EN�G'D��^�X%��W�ئUj�tnc���<l ?��aY9��e7mޒ)�E�Ț�"w]��e�A���0o1+�Rn������|oq�dhU��%��o�ӽ�q�\y��%�c����1��/AUX�5���O��n�3-��M����`'�F��N�����?�X���ϻX9�x69w�-Le���l�f07��r������0�y�L�vS���*������[�S|%F��JG�.!�_D᫐�8��
�j>V���7%��2v���e{hj�����[Tl�zu\A�X]�3��� я����}8����>������}&�-����2vK�$םS�<Fd!F'>�BMDև~�8j��ɽw<h�qn:�ө�PdQ	�獌����W����p�ѰPצ��	�>��P�&�u�~�}Nx�2�#S���I'_�F?<']�Um��d��l#K�'y�쾴:�;/��uc(۪��ؿ��H`J��_�������
�@��7����a�F��������%�Rq}��B���e~q��ۮ`i��ms���6� ��Z��5EjfZ��/�bu��*MN������΃@WK]+}ƭ_Zbt�w�}�\g�^��Wd�l����J�;Oh-`|u�X��}�4�E:Qkl��c�=�M{{@t�Ǳ4Y��"P����� Dރ��z��0x���I۝ٸ&���+��i��j���r��d���9"�GجQ�ǔ�׸$��PI���pi�a*f~���d��e{�����R䇇���f�p΢;�#���[�h��li�%m{Q4����k��!{8$�{��� �sH��ai��h�T�]���N(M��~�JFv}t?)r@ �in�Hog.{�4����;8��TM��9�ί���)�zZ���yPP�U'՛*�}�@��%܈5J�,��8��,��L�(�E�^�ΔW�D0^j���o�N^*,��'�ټ�7uŜү(�m�65LS%ʕ�Pj��SJE>!n�d�à��f9z'n����a�x����
q��v��Z.��25�c����pY�5�t�/O5��@o��:�5�^X��l* 6|V�����X&2����'��b�*�F[y���3=��s�S���7�_��/fL�dU7R�8��z�j3�(1����Tv��Ԅ.?�����ꮌ�4Y[W=�+�%�q��H��>��<1J���^��$k����Rȴ������X2��qC8����x�u�}�{>D`��X�	_M.�Л_�9�>m���l�b ஀2'��R��7�[�7�j\#+�c`���
Hq]���DMG��;��ohh��s��^���&��0�s�9��۽H��jL2!
��V"�=��s&  �61Jm������n ��H��e�v[�����/P�ȶL�7��Qd!9^�s9��Q����|�U����yp��X�JGG�v�i���i7�j;����m���`�3��x';����װ]���Zhӱ�DD=b��X�A;xk�h��st�����E�1�O�z�4��"�/��o���G���B�[���Xx�]�u[h:x�`�x�m�=��Dl�{Y��9hA�����Pq33���k�{�ptoJU;yAV�[�Dj��CP�zy���A_є�~���w�`�����Qd��=9����.��g�Pa�?
��{�_�,�1����kFi����	g��u����Z�K���To�O�� �R�;���Վ�S?2f��NǇW��G�̘�x�=2�w�PQW��;�@2sqR�:���gL��VK�cſ�g��8d$�P{ʲ�e��]W�;���`�$����bPt`:ۗ5ӹBUդyy�F8�ߍ�Efy�"hvv���)�e4�ޕ�7~�oY5)ǋ�oOK$�.���j�l6 ��&	��l�
$�\?�r���h�YkaA�V�r��p>~��$-k, X.sx��Ґ��6Ӳ2%%��C��_D�d��ǤbT��Tz6�B�_�3l[àE�;BD/I8/��I�>�I��$�3c���+7�}*G������Ǿ~�Z�K�ho����ӓ�ߤ��W����`}2���}�\���w;�q�P����	j��k��t~߅6��b�6����:���^¥G��!���l�" �4f����95�,|���������2hA�\ �*�34�7�5��J4Wԗaz�����tU��e���$�MHo�N0�Ɗ�����C�_u�q���[~B2zo?"�-�u9�(d��%��O�E{�<��v��V;�u9%s��G�^!���	\-��x٥c��Il�'���s�E�A�fx��(ۙJ�D�gg��65u�j�g8�]��z�M� oa!27J��!��w�Nw*��8���{���Pf=ߐig�n�D�P�����i�tCJI��ӻ�x��w>s(hV@�8�~���l��Xc�⠢���=��ڹ�3������7����[?KpJ��C<8G�����JnlSH�3�B��% ��k��A{~6�Ҩ���N��>�<����8���,(0{e�1?�0R9�ܨ��R�h�E�H�="�7*��D��r�7hq~�V��=��:�I`%^��ݬ������5�QNwm�z"z�'���z.w��S�]Vܳ�y<��k}}A>T9,��^�P��Ye���(R5��������.�����w�^�@P��z�k��t�-~���q�e7���"���� �g�C&��J�=�X�7r-��_�ǌ�wJ�&7��<,�%�Y�s�Oݠ�Py�d
���\���Kc1j$a;k�4����A�$�MEUO����2��9Ȧ��z�����\^O:CV1��eT\��	����y2Ӊ�m#t�<��$qrn#yfؗC��M��	��!	��G�!#�2��|�i�ķ}���9����U�9M����gRP��Yf����҂;��t��j����A�&z�DkFǅ�,@��s|U&�����E�ͨ`���N����MpH���nB gV�H8|�`�ɱ���h>��ޞ�I?�lc�$�Ê<�O��ɤ ^�>{IҝZ���+c��_7 �����1�ۡͼ��W�����^"���A���6�:J"!>Pjo�/�Cs���vd����~木�{��>�}��b"���rhzw�ѺqR�#�x���jX��M�׼�˭�E���=�T��ڣ��C��c���\��U�����
\�D��W��@" ���7�Ү���яz�/�����7N>��r:nM�*�����5'�\����H#ꕻc�MJ�6}���
���^n����S��ǇJ�=|�K�@H q�kBS'@o�Z%(3e�ix���,�y��V�E1P�g�+ds~N��V<(SW�� b������=�\�t�ͬߢ5S���S��
�~�����MO���dO�0Fz�ޓjV���E��/�3�zm����sHD�@��ޢi�?�/4���]ȼ�ZWף��{:���P����'�4:�7���b��K$9yS�Jr�VqF��u�ȑ��������O�Ő3E�cӼ̆<�[�6e�n� 3�|.]G�T����,���G� v2���J�@���<�U�����AG�;�� �sD}:H��:�x��h�� �)K�w�b�@����k����������]�ʘ�JInx{�'�Ǐ�d�˭?.�G2^�P �S�����Z��p��l�":��+Ǐ�Gd�<�v ]Hr�y��oc��/��uZG�d���t��1�%S%=z�FRo��jݑ'#� �M�oiB���3���	���{3zm)���<��4��𕥸O)Q�����t�T�K�f�i�3d?逾y�D�BtB��ګ~Wz6�>�c�h�HO�����K=J(��+6�� �S��-N����:	�	�\��:�AMց�U����3pz}"Ff���$duH3G�g��9�h��-Ď~+y5�+U�sQ�fw�;���,C��d��K�.��pl��\x��l�ӌ/K�J�'��e`l��pMy�eO��m$��s��D"čk��yq����UFڲ��+�ƄƵ>.�D��~	Nj�0c;F
�孟f���ŴB��+(���]���Ȼ��,��%���Q���2���wAݩ�@#vG���0����R���kn��%�j���0I��(%�l�n�₮��r4��߭����m��=����oU&�U_Z��ݧ	u�O��DK��+���s�P�%_�q��:K7�W3�R����7�Bbi��K����)� y��8�h�} ��\�)ts��3sl0��r�7X<���F8ð�����{D�Sۚ��E�x$ɞ�S�+ -u�G��[�y���q�@���8���%��k�#<��o�z�+sv��X~�#�6l28/�#8��J��2����k�oZ�s�X���,�h��a��qRG��s�{*  ʶ�	�{k�EK�#%h�����O�i-d �C�Jdrp�Ը��EJ�;w�nM�
@�~��X��r�X#�}�����B:��'L��b�˹���3��孢8X�Q�NcҚ�@~��r�;�w��^�	r����ݠ�>q�������ų࢔���0���� �8aaJ[Mm�۾M>x��M_g��b�i���ǎ�aя�̙>�d3�ZF2�VL�n� g�B�����-DFMhk�A _ųY��R��.���Z�JrC}�H���8E"�0u-mU%���9fz5��AϝO�Dα?�#���1G*��E�Ԩ��h} ��\��LH_���!T�h�}�����jw�^��mj�\���IT����7S�0�w��ڢr;���:�)���b8����T��Q(��pֹ-cn��iy�Y\�C��^��B �_�������gy1���hv�'~�[��NV9��ڀ�99��ңy������{/��b
t1����<E��c���O�љ�������0�s�e�����5��9�H=:l$��> zXb�X�
�����>Ѵ�b�d�����yi&��m������.<1ᝁr�s�.�F� e�<'r� ������%=�]��^�}0(xHa԰ J�h���)j �s��V����H�B�n�s��R :*�wd�̰����5 �h��#җk�{2Z���G�=x��{�d��*{n�^eq���	x�V$[�i� ��\�f���.���@��=26�;�r!%�&o}��drd�kށ��y�������p/����8���Φ:!:�� aM�6���rh2���2�=ʹ�ڋ�0��.�2�.�p��~�v��<�~���U&v�Y���?b����7�!),�.���!�~ꐛE���j�+�o:PFҙ"xAޖ�:��9M�ڷ���ﳊw�pyv	dAs�����	g����3+��^b�+�7�Q��G-�?��Ϊ�w�߹i�Z��N�ۇZʼ�e�?�����u��L�|�bV�>�U��"����j�z�0��`��9�������v������5���̬uJ-PZ�$�( �zVPHt��y�K�|,)5��`�k1t�x6t����ƇOA��y�P�P�<�1��V��+�& .�MwFO�ғ;�7�+yO�fM�|�����:|��T}���K�w5�XUl�Eo"�U� @�蘃w���-��r=��W[l5c�
��-���K�m�d>���i(V��'���T;�HN�3O*���6�8t�/3_��+�����������H��T���[ݩ���2���!����;-_$3r�HL��Wr��Tr��d���*�C����̑rVi�.I��}���e�����5�oXZ)��'�3������O��޲�x�y�Sd��}�=��w�}�;�q@�u�� ����#��7�ꯓ��Z�n�����`���~ ���ʠ��^��{�2� x��D�65�	=]��$P�K�2����f���k��&�$'HT�[�}��>Z�����>�,(#�A��Ғ��(ʥr?ʃ���h|��2�M������oH	:_��������lk�i�0�I"��1�yS���$`���s8n<:
?��r���F[ù�m��熻�&�5l�l���ݵ,��0���k�Z%�9�3�0��;�-����<K(���t��z�܀$8�Q����M�
"\
�k����@���V���g�M��Kpp��9�U��C�" ����\�),T�c�acu�$#?�	'�0&扉�є�#%UGUn�$U��y�NE~U�@���A��C�S -84�k�?G�vȂ@� G������'��G�L
�F�v���d�Ă@FYRE�����FK�'o��|NNRP�������X�lGGTg�ҁ��f߹Jx���1䥅O�4�4�6�S�VGީ^�����o��<��z��47ˁ�]VfɸaTw&c䇡��\�i�,%|}�U5�zq�"�%f���{�7�HZk]&�w�4�6�ٌK�̯o#�g��-���'<���8�
�;-|��ede�zR��!q�|V��� �i�N4I8��ot�b�	���v��Jo77JW_EG�D�_��:��H��{Ň�2V��pu{����8�h1 ��a��^�b�?��'[��e���L�y��z�;�O6p+�QҤ��7�z�}���J���A7���W�5V������R�_��^���b������G�P%��֓ϴ�L���1��+:9��Jty�me�[�7{k���&��!ľ�]�jwG��/�@Ŀ&'��&
5w>��,JO 	���?ͬ>��}�O��\��0������Z햂|���K �9��F��c�U��!S���o��xR��v�R��y${АV��'���^��$Du�@��KP�H��<K�3��~0�v��#�/����k�_��s`��5�Ԙn/������J���pf���
h��
�/�_���������-����B��>����T��z��%��Q�Q�:�u���{~����A?��C}�=���c6y�X�*A?���<S�pG�ed��,��A+l�����\O[G��\$���?�b|�4+��E����FJk<��6KQ}Q�Y㴸4�$��'�<#�-�K��p"��#�9����H������ש�i��6E��M�7���auӼ�3��7~��_�	M�5����{p)�*-5���-7�HWOK�7�1�>��0�6"��(����a~X�����+�e3^��¾�V0�i�hQ�p�z�����vgF��Y�<|��Շ+��(7����n]�t�����x�����8�Y3,�����/�*�x��Y7���yB��׮"�^ܠ|��]�dr"���w����vP�(1�"e8��m�ڱA�UG��K�����!m����Wp�oo���H����d�h�`��`�P'��6G��˓]��S#ć���ǎR��jz�9	��E�M��yѦ9��?���C��j�>������ta��^��73��eT��h'\i����v�����S��8v�5�=���	rgav�HwW��_�)x������y�H�ֵ�2ߑ�+Z���݇���Tr�ꚴO:�JcY����g�M�\��UP��:�?�V��E�����9����l��RF^�|W���fI�9I�ڔse��Ή���c��:6$�n�f5�l���l��,�)���(���%'���su�y��7��w*������o.�ΣF�����^����+Nq�CX��L�PI������	t����j�rw���xF����_��������B�im"�����\�yc��oĸ���k�#60�Z�$g��B�⾴;���;������U���Q�o(R� |j�^�O�k�8ˌ6$�5����w�c�k/��W��ނ�+�cH�쉿
̮�����C=��7MI$�]I`��kס������Nf�b��/ЈW��~�]����ƺL*2������7�c
]��c�j�,��d;-e>�͔�ۓ���@f�����4�V��g�I D�'�&Tde��Mx�:��P�[��_���[���h7���|}C���y�#elO��w�l�vT�澽�酴�ua����4�@]��29��in8���x (.Ҕ#V�$9�jF�h5�
SS"G�
ّoO�ற��Xi�#_<]�_}C3c�޼�=��q9���ܔA?�v
�?͗��u�<:�-:5�P���Ĥ�_/z��Z>��"���}�R��9={�f�>�f��ըz!�8�0���D�����Ϻϓ��孶�0��5DH"���K>#ӂU�Q��` %������iW�P��a�g���8�Ɣ{��&��i�#���l���������r[}���+��Ǫ'������.h�)}|Ӣ��I���-��Id&O��R�'�������9Ɲk�:7!>α��݅�m��Cm�~>=�{<� �.kY���)�N�*F�8:��i��_6��1�َ	�
��[����4/U�����l���36ޘ�t�����2�$$���V�qT�ҲZ��p3�^̶��J�w�²ۦ㭶��;�;��R�<z�� W] <�'��"j��Ph��uߏ�4q)��6��n�M�$34���_vy^�y�DŲj-$r�fvk9R�������+,������Z�"�i؍�.����V��?���H��_��n
����= �+7���)m0�z�����Ws+뛿."�$���Z�x^r���ȡcR��v�ǋ6�l?�I�?��ڥܧe^���+�)$Y��vMT�i�A�CW��N�a�6�{U��	;�m�9���Ek��b2���>7���M�mia� ���O�䪍 �Ӷ	��~t;�w�"�֖8���@s'����AZN��x��=�:,����k�H���~��p�ӻ�·�w%�iV�Y)����®Ξ�)M�w�6��wF	���4����]1���<�X���,�}dK3���i���#���o������t15.G�޽�����C�c�Rv[�M��*�5��+����D����G� L�J����궜���ְ/ߤU|����2p�|� ۅ��B-�Xa�~��jƛ�C���o����YU��Y3�A��<[���:U�{$�X�ǥ@�ʟ�D���
���_~�6H�����h'�{#:"�����E�F|�Jb܊�q�L�om}u]C��<����p�$�CG����<W=9N�}t/�5&�ycj�@hi��H�ܽZ� �.U�j��/���KXKv��F��e;�ŴA*a�cA�~$@{�Eb	s���5 !9@�-fff�a�.B �P�9�ϡ����K�yޒ�s�*����9��[��s�17�;���~���u��AP[�v���U���V�T�5���8��>�Zd0
?D�����c�Y�J�cг�=٪�~B�r��7
��\��Ѷh�JQ�<9;)i�O�Q��E^��:m��+Q-D6�D��,*��Y4{bi�E'�4 �	W��qj�(�u�4h���"�����H�ʔ�:pX:�5(�Q���5�T~ӥ��h��U�� ##�'Ť�p���K��n�p��> S�ʁ�y-�lZjN�`�x������߭K��;��Q#B��F�f���]#� Y��U�`T��ӡ�k��q6KȌ';hY������;�]���Je�E��}�r�_huB0?XG���O%�t���Z����~����������l[�h]��[ZE��� a�^�Y�!�v�c��v��m�ܲJ�_�F∐���0�ܣ�w� J/�;�5�D��E ����h����B�6jN�����K��En�C�4�L��bSt5�Wn�ĵV P0#v�t|��+(%��9�>��i�ψ�1B�?�X�o�U���9��ᙤ3!��3��)\���2�s�f|i@�� �i�9>�t�C��VJJ�J�S5���e�r�}����n]��|'+L�.�:�_�n��\�Q14��@������c��̿"y��_w��`�`��	��=��y����{��,�U���I�sZG]-��� ]�!� �E�\i}�NI{:����ϮN~7���TTt49��"�"Ч�������������?�m�@,����)v�FU���b�D�ˆ�mM���9�>c��d/G�ZZ�
o�:'�v��k�R���f��Qh3�NK�Ie�����t��?��&�&OQ�k��aX?��V�Dgh߻�B����;���W�b8:���ɮ!>-�ז�Y���7|���b�mYa%?g�� �$6�
�a�U�a�qS[�<�r����eO
��oI}0U�+���:�9u^���@�%�W����Ӛ}��H�Ȥ��G��/ឮ��S�Ŕ������P�v}˸m�W�{G �S�a��0�M��J�`���w���ԝ��V4�f���d�?�(�y�<[��=m�$��c�g���qy�GX@��˃N*q�םLh��b�N�y��w~\���(ݛ�Vˡ �k����?���$|%�~���`/���"�'��f�)�l� �G5n�r.�PC�����O�Haj[�Ij긍̉�P��t�a��S�H�o=�]+v5�0�%��c�vC���*���I	%�w���a����.<O%�5G�5��=O���Vu'�/!��XD����#��P���%Gl'f9�C��Fk�K�+��q�Kg�.V�LV�?c~��,4g΢ߟ�/�< F˿�26(������iX�F2�ojኦ�[倿	�N6�"m[�is��)���̓�����|����N��P�2����lhU@^{��{��W��z�|�a�\�f��b2F�@ݶ�k�)�y"pW�_��r��flj�ר�g|���F��D`�6ѯ	���.?�O4�*���"�o�+HO�����/>l9�����T ��{?=k��g�P�9���<J)I9✮9tmu����>>��v��6z�q�*�L�A�F�=�MI���K��۩$U���C̆�ola�|�����t:��r�kۃ�n��F��w�w����-�GW7�-��{���.�x	G"IΕ�C)���y=,4�������S�3��s�LK-Ø�����7@%
jWa�A{��|UF���2�"Ye�������5���緹���#2��!ޘY��IF���G����N��E$7�~��d���r�S��_�U�晷���<��(�4�&�~�Q@��9��'6�X/�bbM���J�J�y�Y_7�U�"�a"�߷Y�7ֿm +���\�ѡC�2�������[w�h�������1�Z������-�Aݣ�R���>��4���w��Q2"a�덭^��<u���>V����Q1��{b�\�ISz)�̝\�)Z�$nM����^DqU(䰓���F���U�˗u�ur�"�t�M����=Ğ%+ �LM?ON�Uړф�)��*��3Ρ݋Ҷ�����Cr^m�T��'�V��1h��6 >G[gv@L�Q��J�)������U����s��⟌���4E�u+�t�S��g
��BF��^{�en�}eA�C��S����;�-t���؋���S�

N��R�(�S��<eXi�(��c��?�R�A��O9��Ā
_ ��2� ��=�MH�en������ED�b7�L.����oT�i0@�ޙ��uK�X��5�03s�&$�Z�� n=0�gn'����#~}Q�B�B��W!�/�s��e�(T39��隈#���-��Q�ey�G��6�D�J�b�"9N��ii�]t�����]2�t����&VWY;��0]*�)��}���`s���v�� ܖ�m?r�צ�|�#��hG*�O�fl:8���KSV*1�-�my���o`���	���{(���N���#9f�!I����s�Y�-f��&��崎�
Y�#G�N}�`J���\J��h�P����)����&�����*EĹ����TaDr�0�(md��S�߭^��a����U�_S��|�塀��a��Ƨ�c�|]�.]I��`�����3�=��sv�u �Wݠ��'=S�������BJ�V)��ݟ=�2���_�:�8Vſ���aQ�f���in�;@Zysw��|�cEHS���c��G<�(ܸ�����ﱑ�-�u�1�XD�-[��d��#ۀo���Ƥ?�~Ykg;~�>8u및���>�.9�u���֜K��&uF��+<c�#�v�+�B@�OW�\���q�ٽzz�������ǫ��2���o �_bU��6�*��N�r4̿�g�����j���mF�ZhC��9�7}Ҷ���r�JFE�-x�l�IL�������l���p�b{�q�K���h{�Y��5n�F�����S�Z��Ǽ][�;~�r���3��S���	e��*�!���U������n Lީt�*��>{W�Ζ����e5`.]�P���M��i͋��&����ʟ�]^�k��\�]=[������ *��}x�bTIU\��O���up4N=V��l���l���y!~��S���`�
S^PH7ڢ���/���Ҵi{�DD[%�#,��Уl��t�pI8ߦZ�W��u�B�H雞��.�>Q��o��	�g��`�ՕSVC/���(^��`��6���U�,�U�2p���/L�����p[�ydwx�q���[(�5N�~0��U�!��QV6zllh��<�%�ݰ�Fm�@�5>~�e4#b��@0'0�kS�5��߉MHJ�u&`t?���d���Ȣ@�S s}hn};-����Y��;��L�}���@($^K��b
2�DI�,��T����s�;Dv�w!�Z����09�e^-��� ��d����ª��OK_�TlD!36"V�ʢ
ɠ�lqh�B(����nĒb��7u��������V[]��VX_{���3x2�=��ٲu��פ��� ��Wv:�o�������;V���H������4|�"U���إu�����h��������9畒���Ww���	��v���ZKk'Î�T����oH%�HV�X��f��rq����C!��f�+m/�$��S�rhU�!�O7���A�v��s�j��E��5H�+�K2�˷s��ħO�f����xQ5C9�U���o�u�	U�XC@�KA-�����ꅦV*��HI�1/�؂aKBV�cw�T�����ya ����=x����X+�?�QP}>� "�?�2��G�+��U�5�c���NO`������rh���w@k��E��|Ϋ�wq��s�|K�gɾ�a͒�41�p�fp��i	t*)�K]*䴰k�{�ñܳ��*a���ьд�}7�)WŹ�Y�t�:,ta�ա����9�a�C�%F�G\��6u�����e�#��~)��HN���?��;���iQQD@��(*E�A@:H�"�{�EiJ! �I����z��%�wr���~O|��ٙ�k����Q>�u?4�=��~�5x����#�@[1�I����%��ިw���Q��a{��w��Ds���9����~O��ת�s��<@B��D;���K]��'ғ��]��sN�u
�,�� �\B3�;n�=D^������{�M"�:����*bb���E�,��3v��Yd��x/5?&�w����>;x�~��@ ��l�kTc�j�."g!�frMG���l�(!R8���5�;��BX�zi��~��5@7v&���\�:�nSf
��>���,�j g��Iv1(�C�V�Q�`\M���C��*bmV��NK��\J;�m��|��b�x+x�p,��j�t���f;�Yy�C��{���du���se��1,܀��yʢ��pT�bXH(��ͩ$Ӓ�j��L���,��(�F��1lt��Cd���X�FP#�7 x�����VR3YL��睊��>���RE���K��ژa>�����ƻy�<PM;��0��`	������������d��,���.��t��j���n�T�{��ٙ8Ǉω��D�Ұ��4}�MW��;#��]o��-�e����rv~�$̜m�@��hְ�(�?J�+�^��A/�J�X=��]u�d�G�/�95���&q���1�����������,-������VA��2��)�&x�r
dJ��ccr�9�+U[�����f3_��"��ֿ�4���4�N���T�om�����s�6���_�YH^g�AE����tP��<�@�k�.�a7�)� ������Fq5`dTˑN%�B<B��|أe��5IJ|I����_?�Pp�F�y6+�(��f�v�UZ@���hkY�P�)���`�J��
��<ܞIQ}]�G?:����;��ń�v27)K��U�����Y쏛�|
�ޭV�o��C�ieM��;(�dp\��K��!y�����p�@l��x��Rk��.���o���ƶ,���;�?�y��\/�nk�7��o2��m>��.>�e. �W�&$��N*n~��؍��\Б���
۞�=��d���>%�!�e�)�i���z���Z��6=>���U��C,a�8vVj�ȼ���vs'#�L� �ڡ�\�X�j�����W�UrG��f4�]A60�v8V��m7�'h�G��n��3(�@T�]���Xy�>��o}He��V�J�DuE��������~��4F:0���58��.U���@�N6S?�<���/��BW�ٿ�?vA���"^4C��ؚAF�@�G�t)oe�������M>�cN�T���$I<S��-@ի~®4h��-�.�AP_}b�%�3��f-!N�v8mv�֠ �޼���
-֥����ܦ���/�q;O�'��+�<q�`m�E��H������	�3J3��iBȤ�ڐ��.v�s>��	�Փ>TC8Vɲ��9�S|w�P-˵+v�Z�>H�����(�#T�O�,�l��YL�o�:-3W�-�ԗ����n[�|��k�P�P}��Ebvp����}���^��"����ijg���	nI=mPU��_=���j�é�Q��A�s��X�Nc����Z$�'��{(��E��([^�`��I����O��k�j�hN�j�A	F-�7I��u!�m�מoo�:����i��E�<��=mùS�f,��D�~��m�fOb	��.@lτ`���Ğ�'���mU��Q�����l�� �haQ��j������]ϵ���a�;��dZ�A����]bV���t\�(j�ą���ֲU!���7�kYG-�����]��)/Mn�?��=}�۫ߺ��h�7zʻ#۩Cq�7�Đ��wB�!2��Ƿ��([>�˛^������PliV��{hL_��9�BAtꞒ�6-*!ѵ&�OU<D�E\����t��XfXT�/�_S�1�H^\�9��t�y:{=*�M~�c�Z��N��:x�=���ɑ~H�<���v��:ӡ�܄��K��Ro_����
��9C��"�r�摀�b�i2���J��=����ڐژ�$�Z������<�M�7���kX7�?�MD5�Ф����I���H�kY�l�-|����* ��[��V��StV�܁{Z�]q���s���A���Q��I	���Ē����{�`��ﺖ�|�ꚞ����p��Ik�n����V��
�B�/�Α��Ro����_8wm �)�~��S��Y��_M�F+! �������>ȷ�����o��.�7����21��@t�۞����փuԞ2̷���rt�|�����5��G`��Cv���>�aO���r��~���<�mޕÍ�^��"��:�u�;��'�W:���ȶ���%ۇ$*\��O�80�{?����T����0tL�������-�Xk���"e���I�ۅ��&sQ*�i>�����H˗��TzE���Aun�[i�:�y_z�3j��P.��ߗ� ��y���n�{�a�Ҿs��@h�3| "��P외nv%x�c�Y���ԔV�����'�@.o)��xck�2�������&�}��ƾqC�Az_n�{@�n�n)N�*��na?�\,����?s����1Z�zaa���w�j��c�ގn֊��FDF�XΉ#�p~�#�n߭޼��,���v������	~90-%Rx1�����J2D�k��J2WH��\xհ���j���d��lgk��ں�y�]�k������� ��V(~�]ي<<vLH�k�Δ}!�7nɑ�����QP�ؒ���@{v�]Jz��-�T�qIUU�h�/�z>�ps��=��C5��seE������H��5��j�j�
m�1w��O@�M|��	�tq����{��^D� =���D��_�W����j`�:)�v�Z~��>l#���ٖe���kOeS��Ś���;N�9���&�Y�;yFz���a���9�Y*�܁�mmt!�3��;�ܠbz?t��.h�?uv:��^�m3�=u%�:HUUQ���F�5>>�y���KKK+����ԬBY̡�S�ϩ�~!=nȵ>��0������lV/�Ձ9��n�<�U���I�v��ͺ���6w��|l�ڠ�6Ҍ(45J�M�f���� jD�˃sX/}�:K�$ٞe����7M~�u݋(:D]�3'�+uZ�?r���Ҵ$Ae8����<�Uٷ��c]��nW�e���upL�U�d�t�u�2E�)C�hS���� ��k��Ʒ^f:�|,���&6��Y�:�x�m����ߡ���Kp	T�!���L�����@4'8ӿ-�6��q����?�5'�)q��"�|�07M/�\�/��,���6DYU�Xn�s[�_���W�����0��^��m�n1W�&��0��ݠ�� �7�|fKp�c򷜽��8z|�^r��ZL �ӿZa~�5��|�����r�}YL�v~�#����o�Y{�0���R�`�ؕW)K��ʉ��~����N�QJ��q֮B���]��J\K?��U1oy1W�V!�w�����V�ިϔ�����}�v�I�q.�Ue�Z�bj"׺G� P����(E\c�@�U�R;=��?T���4]��k��c�G*���|ݟ@JKO����[D��Z��.*r?�;Վ$��	Ƣ��{�QC81Y1��s�R�:����o׻E�6�'���6�����;S��ވ�n����&�DWV)��:{d�!��,��`��+��< �ĳO�G�9������B���	�2��Z������y~��hq]2�Te*�ku�������t�\�\/��#��C�5��w�|�	*���$���@�t�A�ۤ�a�so��V>��w�$��,�-kЯ7��	i'P.�c�K6����,�>��绯�W9���T&����@y&���Bɻ�����oR�01���j� �2�����������ASR�Y(�)�7��Ҥ_�3^!�Oy�_�s��վi�WG�s�V�aE=9-,��n��{�}4B��������>Z�}U�oP�ؙ����})&bAmc�%��� @���G	�ck/Wy|ד �7�[>�ҹ�/f�.h殭��M\���AE���O=Z�@�v����A�$Pr��?�w2���̑PR�i}�1`ŖwZ'�|>m�Fy ���	�Ϊ�_H�)Fi-ށɢ|%��ο��E^9e�{�2/7�gW3`��p�aX0�+��T���������\)�0���'hS�%�_8��
�]M��Wb�W�EȠ�����s*�1^ݤ�9�m����~�A�t���FfIj/B.Q믍�"\�#ּ��.�/T�r��3 �N�e#��uD�k`��_�u5o.�YiĘ�7UW�s5�o��`<o�s+�b�)��T1K���O��`��XJ�'��C�Zq��h�
�0�{�_�w%��r����N<��3�zy��#�j�vJ��r���׾�/��\yֺ������ĭg�@�]J��C"�u8���k�=�k>J���GK����,g���7⁲Ω4ׇZ3J+5�6K�n�?�B��/�sһ�.��i���rRn�m��ݝ�x)5p�� �D)j}�"�&������m�
q@]Q�v n�wK���	����>����H�2dk��qf��<.�pIDQ�K���6�d��~��!��n�+o�Xr�g�9�Ü��	��؝�?ޡ�����9L�n)β.���xHR=5�������K���n��Dz.M��zO��=����&O�y���I'��hM�z��	���D9;�桘�JW�>u�а�;QK�����K�e�g���%�63��,���k�	�������"uDAjZ����g� ��B��|��D?2O�Fk�R�9��Q�o��{H��BK:�V�3*�s�mZ��uH��/N�7���0Nl���o���x��3�)��%�~nO��\�|p(����_���33��.f@'`�v��	������ <u��`R��S1�|S�֜�z�|����Z��%���t��L|W�Ǡ_53l?��КTr�8j�;T�=���y�pA'���1H�����H���/ @^+�' �+7;Da����pP;�CA~���v�^���&�{�[�����e10���L��o�IE��h�+���x��HvW���2��,���ȍ(P�k˼��q��}�Ǘ����.4�:ռK_�2�<^�7�<	|��k��_���,i��kp��:�
��+r3IL�2r5��>���f����Z(����A��(��8
���&�E��E@j��80	id�[�;�R��w7�9-�h�3�_��N���y��zG��!>��s��8��qo���/��>�.(7�4�B(·b6��w�,���� C���������NO�r��إ܆��J@đT�˖ַ�cee�6��Aam$�]z�G�#�R1��ല�2o璈�T��;]�4Ì��ױ��^��Pp��i�;%J��T-�ԏ�\�hd�-�Ϳ�ݵ�W�$�U���B�P�����L��RY
;J=�K� ���~T����k��J-��n�|?v�Nʸ�	}	F=W��F�4�' ��Ϧ�q�.:����ۮr������ɷ�,��lOVB�d��i5W��ֶ�6�yA�ŗ��d_!܈���棻�eX�����N���$�<0սZZeq� ���_3n���ߜ{~P�I�V�\��g �|Q�^���r~��78W}X���Ħ�*h� ���b��D	����~l�~&Ω��]�aL����4Z(���q�;���_��5+A��ψ���j3��R^��e�:��ts=���b�;����܀�'�jV�p���s8_Q�_p�z�&�>M�j7���)�~����@f�Ɍ)�1A��6ۀ7(�BOZ�e�_) �������`O%Ш���=��#w��f��w$'�'>Z[l�5�4��7��� �ljܥ!�5�D}ꚺ�+�o�O�@3��լl�������k7�<;_KY�</FoU<^�ov��i�����",��$��EY�_j�Qu�Cs��cm�*M��7����B(�V�����^��Ǜ��/��jg�GY����pr�k`Φ�rµ�ե�K��Ш�M����+��r֑l��iy���Z�v�֨�P7�T��f �F���&|�^��C�JLA��a@7�CdF�~ucU�H8�A��7��L��J��v�|��q5��ۣgסD�H�R���r,�<�����9����N+�;����6�z~�C�d��2؀�֮t��&	���C��*p�FM9�{�i8�o�5Z��N��~0Kҹ&:h�4�9�'�Թn���,�f�� Ĉuq|����Ņ�"�]���p�j����5�M�����'ٛ�L\�R���������;���ٝ�t"lGu�Z28B$r�e�w������O��k�)�a�=�!#����s�m���������3_�+3MƠ5��a0�u���d��?����9ݪ�}ݽ3�DN��"9� �N�s����Y��ve��;#�y���D��t
�f�-�����X�!�"\�a��6��?TC���N?���t���P�>��@jé����㏪�gO���6�U�4��N�m������kGW3u�Y�@U~��سZ����_J��+�/���%ḹ��|NraS�u(?7�b�`F)~?O*v����thg�?�Y'§�|՞uD^�~�/-�M��4b�q|�N \V��zٓU� ���}��s\��M��ΗW��i���E.���cF��b&��Ă6�	�@6�J:d%Vr�$�A
��(�u�h1]�>������X{�����/D��&��8	�A���Yf	[����YV�$���ÞNaq����G1o?��){/�kxe�\�kt�J��"m�-����>>r��O��3>����_lt��r$�{���5q���*���6�����=�|��ɵP�rm�a�@1���\,_s�pr��L�e�����'����d���t��Yl:��\�s7�j�x�.��|{a�zO*��B1H��� ����g�V�������D�@����r���S��H�u�oI>�U;Jӹ��~>	����.�5@�=Ó�\�(�K�(kN��"N}���,�v"�kqI*eHP*ih�N��M/� 7`��r�.�*��Ҩ���O~��*J>�4�ҞNs7���证]�S7H��Xi��5�;PKz�˛��eڿ����46k`�|I������39-�Vs<��'�����@l���l�v�x�P�����=4������Aj��m�<��p�|��+���+�П� ���g����	X����u)Z[Q�[�
��*��s��!u�w[��rE�A*�4��b��jiSc�KEU@v� �z{�0�����AY���B�5�h�"��ݟ���Cm�
Q
�p�O�iИ�T���gy��K_�p&��uM�
hu#D|6�@��(�k �����YWy�/�Pߖm<.᯽��J��@�sW�\��֨[�,<+�^����DHZ�?z�F���CԠ��#��jo��=�������;#&��i��j6�0[�u�M��!���J8����y�?^x�M������<jF��׸�1E����`wx��Ԍ��?��Iy�^�A�8�>���Q�ʷ��\9ۃ_qϽ�oSRN��wv�����Zm�bpi�����M3��"a_eMv��H ���KE׿�oT��E�@�3�?R��a��dS�^��F>�ɻ��ܖ]Kw�*RV�a�f���x�q��W�a��.c��9�����0�!G��wf�׸qo��-�S��-5F�R�4����ԯ�)f�|ڻ��<͘ ^u�k�<�8���:���57����D<sY��J��-B>��h7��{�Y�=���Ȟ*=ٵ�xߍ�sSc�T8ǸS�px� $����?n��X� �� E0���B��2k��<�j�a� ����7�R���ox\����E�I����<w��j�8J0fZ5��Ӂ�ۮ���_Jj^�^q�a��b�t���������{7�����H""ɩ�q|mae�\Y|������kt�ĉ]G'/=AY�u�5-�c �3N�9��&U��(��=�#��xA�6:}���?�Ah���,Jb̠3���1�EcI����ɤ�J�U0as�&�e�.��Lp$h9��Qz"u$(:p�nh�ĵ/ �~]sR�������'��r�!{�w�[��gQ��p�i͛i*��ߏ�-]��k�U���6�.&�����\�1t�iY@�B^&�������%"�k��ǈ.���XI���3�%9;i�X�H���7ϴ�lt�0�}E���������tߥ'��wn���oY�[�������C���/a�o2n爲~�M���2=7�<��"��g-��-}"6;�J�t�W'��Y���wr%�	NL�t���t8 n�t܎���t|��|�������q^���B* ��:�~O�X��$�y��v&�(%�X�)g��zC�r��脊����'.�'����ݟ�%R	pٻs��pf�js	%Ɉ�a㹯A��,�HG��!�qr8~R�W��8k{���Rem	pѐ,����KO����B�]W;	���|#�u�:l-S���+����;��=�>�Hj�)5��R�8��+�K'^�N���k�����f_���na:܎�Hb`tD���0��$$47^�Ha�;�������t���3$�(�y��˻X����X�~��2�7:�޼N��f�=wDH�9��`��Ǥ�y\X��luMb�:ɘ��������V�Z���t���x�'����N`�W�e�f�|h���I�����/kY���c������x*bz��b���^��[���>8ȍ��2�1,��eG��99]+�/,�X����R�W���g��)j��C/-�-u�`jw/e6YQc޲nR˔�A��=��f�(��s�Ǖ�H��N3�f��11{��EDS�T�~�wK��|������� ]�^��g���mx�������V�e���$�`��D���7|:�a�ъ~}�T*f��e�2J�Zr��U����~�]yE�3�tb�
���($�����Zj�
�L4���ؖ��COu�Z��TV]! �'U	x_cЗ���w������2��3���H_�����ҡ��"��t�2�>F&�}6`�����-���U֋Sc{5\�z�n��+*4;�'Y$�>��ŵ�:d>W��+�p�}&�N���QX:X�ט�]Ձ*����S��_��/�)1l����が�i9~�Hi�����tͰCP���$]�P������`�CZ�F,�����`w�P�}��kJe%
puK�NÕ+'��x��UBw��z!=�DiM��I��Z{lk/�f�|_v}l���v�B�1Cf*8oL�PR��1�U��Q�P��vU��?.غlZ*����Rg��s�H�k��VR����}T��C��y�7P��\�:�l����ϻ8n�D��ߪzvj2@��q�p����gwJ*��u�;���K�fG�#��_��X���{��.��w��M(�����N�hTz�3m���+�
��cR�Jz��LpYvӄ6���[*%�D㤋�t�G��㲵U@�zQ��Sp�M���Uu�&�����;�
����Q^� ��V�s��gg�ȳ���'�o���oFR�:��sE�ql�i��@a��1��#��g��ٚ���}�{mh*fuZ7�C������l$��>똖�^\��=��*���nx|1}a��V�}�?���e�/�0Ҡہ�M_�:���"' Ȱ7u�Yt��  ��w;��w%5J�6#�G�x�Ǐ�����x������[f��,~|\����8RC^+��2u�k{Y�P9rd���R�WM�nX�ʂ�ė���.�!����Og�Շ|�
��ᣧ����/��s�L���&'K�jf�tqo�u��\� &0�q���*��c��4�=��V�>9�{� �y���*]����7<U���'W[hʅ�je�^:�(���*�Ũ���������`������\����
�c5��f�\8�x&�_Qe�[���%����v�C)z@��r��K\�w�$�ҋ��Q�Fp�U���Z`�}��&��%�ԁ���Gu}	W�ʢ<�b=˖��(��_�|��;�#��a�m����K�W�\M�q�2�d�s��
6΃�<�ʹ�3�5|��0���ER���&���Y����!��1Z����i���i��E�}�Ŗ]�����Z���ڐIDs�	���.i�Qb'�������yy�(�13݅^m��y�{��n2��,�eb�Ҿ�bg|���g>����tk���/�(��֐ȅ��s@g9qwh�k��?-6�W:>v��Qo����0f*��jq{��Y�fi��H��N��j���sɆ�-�C��'\�P��@[���"tyq�ş��	#�o7Ri,!�YbY燇�g;�1BzYl�6{���4�����î]'ݳZJ�͓��t��ڿ�ld�[D��X�5J
��
aw��2Yv��,xw���H���s�Ƶo��>xq&�k?ꙇ]2�~̫���g���d��Ws,�x�i�
��UK̩�8��P\��_����!b�gj9�����?�5��"��/�ܚA��L��s�p��!�ζ����	�׬��n�IV��^��r�M㟤��e�뙩E�3��ďQe�Wx��H� ̣��׬n��H��	�=�\J�(�y�̟����\a#f���s��k'�2D���W�^���2eλ	%�>MQf@^]]�v��1�|���'�B,ԇomuE���R��[�s��DSo����ꅡ�㜁V}��5{O���ᢺ�H�d�Q�YW���M�vX�rm�q��t��[z{�x�^��K]���<ɰ�`�O�Roa}:��^�z�8������_�0���c�V.Jv���z������q���"-���o�����D��)�׶?n� �����H��%ä\!�.J�qNH���[��|�C3�Rvg9&��S�,�$rr0�����$kÙ3 v��i�f�m����Ӽ����7�2q��/0&��4���ڏ�}�q'8[G�ܑ�����ސ�b������n}�׵��Y#4�:L�/�n����!�y�Y|X�:�tDW��]n�.w�I�MsN�f����9W��3d1l�z�d0-6L�����?�k6>�{B��iێ�vƸU�:]�؈uC��q��+�A��]# �����U�Pa��4�l5xH� KG�XK�)��}�H��5<2�H���R��*F��e�k��t�.�:;�kWf���|���?
O���I:��p��bc�,��q�i	N����LGEf6v������Y���Y���N�d�����;	uRۂߴ� ��uS��Y�T;ՅQ%�~����J������O)��n�h1��8��kt$������������o�Ͼ�G���� �Xb�r���z~���;�1�fv�uתE�)��@�*�Q`�9Fo r�=ؐ;�I;ʛe�y>�p��*�$���f�����s�s$���N{�I{��F��8��$��}T�̥G�A ��2�.�,	?�a񆁟Be�����@�s���$��M�̻k��kT7YaC����[�WR�I[�DM�1V�s��5X$��a���C��ތ��=Ic]�f ��"���J]�W��{(����=uvh�c�g��;6ti^9���I�hZ�3@�9G���P����"��~ �5��#	p�J�o
��և�����S��e"��(<�cH��#���\�;��y�YJ�]����]�����{gb�/oi�F�Ƨd���ai�� �$s�2&wZ�-:�_[���=��	�>���P�B��Ѝ��̔Nt&�[���-�_��Z���,�=E�v��u^��=�%�:�d�韶x��C��x�@�����G�����Qi�S�ȸ�=���������vژ��,�X�$�c�˱R?G�F��q��/z2�#[��Y����}�ݺ��g�}v{�9��^wR/�T?�����Ǫ���� ;[019�x0*P��W��{��M;�`+U a�TjW]9��Ƙ�w7�ņ����Ybi+�T1*/PB�������W��B7<.�������k��)G���|�Ԁ�*�=@�� �0~}���{#i`��]�pG^�Q� ��2����Gҗ��M:M��XO��C�8ֶX� a�&�~�`��9�"���}�MV�?X�R��!3���M�V�ڨ��ӂ*���'�*�1P�KS��1	��q+J�`�6��u��& b(��3��՜I���\�c�Pp�����]�������Q=����{"}�-&�xm��MEO|f�w3l�ഥ�Lz3[�>M^9�,V�Y,�O�i3�u��q޳��I�A�f,�W�������?P���$��{|���m���P}B.���J��~��F�`�H���X��9�@i�ǻI� �E}z
g���	�٦O��$�a�Gh��p���s.����ÓSS�0���j����%�q]BgzFjjo]��@�`�'��}�vFuC9Eߞ�S^�����D��e�~'W dBM^+G�'�D��N4L'�Ċ�R9�M��4�ӝg����5@� u`U{��f��u�?UI����e�4`O�p;35��-@�L�?��y��\
,J��n��Ihע[�ϹOlV#��+�@�LZ�� �����u�T���I�/4���lj��3;Y�}������|r���"B8H#kte&�&�c�1m��ݘ���TUp��YSS�rm�m�y�G��� �!`8�<1`R˝(f�L�tġ^�g�Vh�����ܬ���p)��ymWkd�4D{��~!p����d�7��.�Ms�)��[����1�����Sj,�y�����M/��Ʌ�RP7��pq1��Y�?�����^BQ"'��Rh��O��>M��.W`穴C�������"��_�`>(&!�-V�L�{Ψ���֑���\5��O���n8Wޤ��㹢���eD��R��Ǜ�-��i:: �$�i����:�c�IU���.�ޗ45��+U]Tz��c�/E#���%����
QGe07L����� �Nn�a[[�h��w����0�8
ȇ��ok^j�����T�h�����U4?]�`��{�	�����]�0����~U<(��؈���~�����s�����-@�[�5�%�UI@j���S9����ۥ��q`�Z����y����m^?+\�6����s^O��yj-�ט��I>��m�(3��e<���LPz%,�7ϲnC[J�fW�c���0�a��S��v��6�(O���yz-�a�����Y��`A�>�U{^�:c�m�?�e�V�����5R�d��zǓ�j..v���=������'��y�P�f�XWs��:�9k��:��_8yc�Y֟1�{�Gj��ʊ�}K]�sl,� ��A��� ��6�����O���VWi�r^����jO��J�ĺ���2×���?��NQ�����5w;`)��:״�X��
��\y8e�ݿ8�5d���U�{B�śe$�!uu�����r{�oaG}(���\�7rx���8櫵ӣ������| `�C���9iHrM�κ�՛r[�-�9��!Oxz��ln�a�k,��ewA�ϒ�w��-'u�Nke�S:�1&�}���7���:eިX&���>��[���������,�FQ�*��խ|"�����!n���y9�xS���H[���I�kah�ⶮ������o��+�^&[�-Y�6�m�6O/�<�g��F�~�,�=��O�#�#ܗ���x��������i��8g���t�=�&��B�عEQ�Z�yS`�g���޹Q�ص>LK�e8i6,ʦB�K���~k���W�:�GO�ӓ��]W��AK�
.o�]�˅�Z&������A�!�c�_�I����PS<��}T��q�h����Q�.N��Ӑ�r�w�xY�c~�l����!�Q">J�:����RmVy��N�b��-<�ƮAIP�����~NT\�a0���Ӱ�|֮��
��6jc��jXΫu��,ˎ�7=� ��	�+��op9�֋X��zx�T%�:]��<�Sy��⛖SY�zT�c7��tSLW�B��t����mP��1��f�dMu�1�G��YHN��a�3�-���K޴o]��P's��6gm5���ٞ�Q�JJ|���v�7�� uj��WІM`��D�7�R��+2S�/�]�B���Ⴢ����jt��s��<�"�+JQ�4��-j����*���8��yӗd�?Kl�M.x�
!��ڿQ����HT�v��r3�Χå9�5�<��0�T�D4J̢*R� �򇳛F>�]��;���C�F_~�0~��Og��#�
��W�+����gk�2�>~�`����KhhW4��RM�|�����ݴ�lo�2��B$p�D����@|nFU��&ډe=�<���Lc/|'v� U�]q�l)�����
i;=�o�^}+���I��I�3�����;x4C�1!9k������m�Q�n�����- �&�9{���IE2�_�ȨX,p�~v�����PS�����Ԫ0�(.�= WQ�/���#���7yٍ��md��������'<2�= �y���B�ߪ�.yw҉֖�	*���������(�ځ/%?�\�;Q�p�L�����I�~g�QaL̛Ve�o?m`^�%�.�ж��w�LM惱 ��R��N���hJ
2��dA��x)������i�R�n!zۻ�ۋzu#��V� ���wD�]#����ė��o~�tٌ��=.����BoD���b (�l��.7��NT��1�Z'�35.��sd���X^;���t�=^�-B�VI8���Mݮ��)�Y��_za��}lf�C#���YY����I�ƒO8�yC��\�����'o÷S�H[C|�̐OIJ�z&p	�g��^�_#����%���|m��Ȁܬ��w?�ٞ�h��Y� ����$�����̉�:�T��*�zb��4(���ܯF������ �fb��_�z~�>����2Y%�Q>�E{[K(Y�1css���G��g�D]�B?�P�������a�����*U}��U臥Y!7�����!NlsI'����ՒYU޺�2w�:D�[F:Ո_&E�|����q�����b)�K�)O8�/��p8�m��ډ��~5N��_^��?�o��������2$�.�+���mfI��[���6_�tՑY�O7z����\���]'Lr�D�\Bw0��}�;#2x�<�%I/���1jA�Ƴ���赹j������<l�7Wh&���e�ʽ���i���/]I3��F�7TQ-? ����@�!��p�!���Zs�Ԣ= ����[���A~:��)O
l�j }'��S�#�t9I~��GL}ɂ���v��-�}����w>�B{��K���??����	�O�dk�2��	_��9�UvOn�vN��/��a��6�ׂX���z����$�FԂڙ����s�u1��$�f��6�)�L`�5Z�L�aT�����Yf=4緜���Z�l� ��I�!hc�} ቻ���DU�I�섄�򚣺 ~��c#��b�C�k�7�� ѨJ����RUI�0����#�C��K���>,{<��~��*9��<3�ފ���=1�����
`N&c�FA��AYL�=!�}�� S����L���|L�FD�Єs��9v���&�����{tT�lW�z��G�31�v�Oמ����@OW�� %! �j�#�܏�����c#I�#X1�K�
�Ա�6{��`+�qb���݈H����:�ƾX#%Ʈ�Z�� �$M[5�x��ܳ�G&}��8Qh�Ë����Ғ��i�(u�qΙ�1�Ɠ'M��(qU�Jj���� �1"���B��o�U/!3�	d2�'<�Z'Z��`�ǡ��=q�I�ٳK�e5��g� �)Y�_js��:Z��?~_F�5ʣ�A%�1ȹ�f�\$!F�d_���v�c����J����^{*�s�3��jD�~E�a+:�j��q�(IS�
��94!*�UKk�5n��o�y���+;��j����2i6�دl[�`��E���bA"j#��'�2����)�K,�aL���nF��f�Ҍ���I^�[�X��v·�j,�L��=���|��n���� �}���Cc����gl=>i�%���zN٬��ޮ����,�rz�K�2UI_��n��$GN&���V�+�>fwGٻ@��Tҥ� Dִ��q���ẖl&��Ju�L��4*�֔��"��zc�ֱ�\���qdX���DƷ����sǲ���bx,2�3��x�{�EZ���~�g��?ۇ��_ �ux�O�{[�Q	V�d ��Kx,�j�YVjXĎ�e�N����[�,eGqm�P5��i�[�i5s�F��o%.��v�3f��Z�M��H��y�v�x���k�NxUF�]ĬH�aҦ��3��$��Iό&j����4���=h�A6Z�X��>k{ �?����|'a$�]���ƭ�_Y���4�|ɟ�RH5��ykVך��g����wc^W�������&��Bء�p����Ǜ�D�O��+j�����][^͍^�S�C�����L)o�FXY�n�W��b4k�}�n��+���"~q�WdW����:K]�ֈ-%OS�2G�9�X����ť)Os\�XA�t>����f��_{ �C���]��՞�]����,� GC��^�&� g�9��3#�
r���X��pK�W���m�4�[�/�a��!BW�����c�O���[d�&��-r��d笓��6�X�"ؗ����1.W�DD_��E� �0O� Σ�����jB���=e��2����P5�
L31���eRw�������W��z�j���P�紈�\�g��:7,.X�����z��@6����t��b��Ӣ�jt:��vZ�(:c�=�%��.EmU�גFKCQ��Z#�� ��-�$�䋙���|�&����s���s�s�s=�rMMV������=���]Ad�x�]�Y�s>B��v������5����B�@2
��HPr2>�c�\�O��B:�7�i㯼�M�oǰ�;y�Ȧ��lܹE����I�V��a���у��'ݤiz~�Y�Rի�{Ҍ" �pdq�ɕ�X-�=�5_�`��`Є1�6z�'tWB�b�P�0��i����|r��ҙ+�)���#�N�2���~-���9����!��5�8�
�3��D�D��s�(��A�Ӷ����x����s��e&�
�3fH��/�h͐�0��Z$�2K�F��7���yݏ0?��s�K��r	7	6{���j��n���g\x��n�a8}����|/+(�a���@����LB�$6�ȠJ۴����B;β�)�|�6]u�"�^�|���@�L���GP�9�)�]����d�m�6��>-�q���#�e�x�*k�Z�-�eo�kj8Q��fi�L ���&�u@}�p�2(����dףC�Cu���A����_���ێ���~îY�xY�R����x���~�q��`u�]�}.j��&���֡��c,�Nt��i�K���c1��N������7M}��!�cvq&{�j��8�����k��� �a����B�ש�Ӎ��k��k�2L�=��;��A��fԯ���� �}�/~���D�#6�hXH�SC�u�/o���m�����"����F�eb�|jK�����P:�Q�~vq�?#}�Ipܨ�H����+|���;�5�5�=������ʳt�=;l����5�� �dx��I�I���Sb1�5�b,����B�C	&�Ze������b�*�:��i�}���KL�OZ�	D�p��)��
B���̼M�EndCzf�C6*��EuMy.&�HU�iX8w��DHJIA"7���R�3}�t�\]���>&<����t\D#�H���{�ą���L�Y�`�F����r��.u�~�;wxe�I�ͦ�?�ҡ��vO��"���0��7I�0�^[R�KG�`���B����N�T�_��p�xN���~�^N��w��x��F�a�P�6�ؙ���Ga��ME���/x)I.}W�]@�b�Ak9��X��R�?�h��Ĺ���
?<9�%G��*��S?F�Jl�SӍV.��lfg����F���J	<�����A=[�4#�)|c��n�I�S҇y��r��!���X~�Ʌ�#v���mLB�|�/#V�T*�!��g.C�@��*�����rK@� ސoX�h+?Eic�����k���e�#�c�o�Ƴ�~�Nl,Ix4�}0�w\xϣ%����T�0r�o��y�"t���#�v/P��B�j�r��W��{ .H݄fG�׼1��b�M�籽���y�@�m8!�����$x9����c�M�Y�>��Q��bR���id7��__Ic�1����99.g>�{	��.��\��8�U����5��Z�^��Lj�D��mX��
���VQ*%{��c�����eY�((=ZL8�J��i�DF������_�-��U6
��j�~O���n3��3�vI�-��%P�L�Ѐ8�gcR�7�̄n�t��.�b_g��m�N�U�u�c�b�"ʷ��<x�x��cFM-��=��J��V�`,3&�=�C��)�;UG���葢z�%kϐγ	��"4c��]�/�c̙	�ZT�Un�{�E��K������a�UYX�$;�b-� �27"g»�O��8"S�Ҩv���N�ڦi�J��k̷�C�A���r� �u9�MRg�a����N�%��Ιe)�����N��~�i�K�#��ƌ �U����tn��'UO8�ũ�Bo��>ء4����\�|�s{Vʡ�o�X}y��H��{��[k�E���<�;d�^�;G���~�$��ل�4Erq����|���&ެ�^��p����)0��Oߎfj�����|T���ׅ�ZF8v���Æ�KsC��6�["���w}r��oZAr(�uÈ�����+,�ştV�/��k�Ɓ��;�:��N l����-,%�Џ	�B��!K����'Y�[�$q)����������N�ax���`��V6�]�gğ̮�dg:Wr�<��ȡ�F��T���FX�W�������i|$���s,Mr�o�R��ho�>�[��G��^��Q�/MɊP�����;q�z����j`c�V^��]!��^�{<o ��q��1o�`^j'�Z�b�������{�Y�_�$[����˶pV��L�:#!�o�32�1G�형G��y�Aޏ�M���Y�8 ��6�Ȅ�|X)�ND	6���P�h��4�Ž����֗�^�� Yɹ��y� �0Mp&h��u�-/�׮�� ɍGY�aW.�?^h��f�i��Qf�T���!!�<�H��e�/�1`�D�kT[&�p��C����":O�@�O�4X����P8��^�0a�K�C`�!7�5����a��~S#���Sw?����+�7�t�+t��^mI=k�I��Pݧ���K�J���˞�9�S�;�if5��8U�*J�vG������#��FڹQ�cO2��<�^Ź�14T�ܤ��x��A���x��J�"��s�]"��&�j��F^�W�ugX�h�ybGp��o��}~eҦ?ٶ��&���%����͸����>�䭾�8���5�^��7j�#}�ztt�Hu9�9�����1Ĉ�w�(�:	�������G��9�ou�_��N4a�ő�Y�������R%�C�� }�_&�R�����T����v/�S}\!?��&���o� ^�I��QfcW�c��r��3*��j�aBwJ ;
��N� ~��:W��ZZ&T�%w}������ P}��2�� �{5���{�7vSL|*�����	�ϭ^����}�zrρ��8�%+{��:�wj�pʜ-Sf��*�8lZǚe�3�����(�yc�u|^���R��A��i�Ѐgʀ" ��-����3eI��1��:��M��À��]��{�"�/�4ծ���o��N�����ih	���-d�ѸU�9\��cUd�����=����8�31���K)&ĥ���mtD�/�]w���L�Tn�!����z��{���6mδ�:��
���ˬ���A��~C��	��ڲ�\b~���umGCv}k�)4�K�R8(lsP���zTsnZ�MP�����o�,%$Ke����Bo/��Pj�V%��o�4�u�Me�ʨ ��6=��!���zԊ|�@)�j���xf�^Gf�E�s1����-�{)k��J����3�}ᐱ���M�Z@k�^�s�Z��	N�A'�Z��D�e�#:"D IG�����tSF�|&O���.�
F��ۺ�Y��:�#[C	�7压m�-���;F5��r;@�f�Tl���{eR����̇�bN��/�u��b7��C ��sZ7�Q�_{3��|!�g��m}�
��M� ��[yy��f�B�`[%�o�]קŇN�$�L(p�-�(^|./���{.ۧ�8ӀB��D��2_�)~i��M�2��y��D��x�O)P��I�2�z
:��qKԈ�W+���J ��S�d�>��c���D����#�PұY�q��-m-���.�!���I�1��{�/�,�֗3z�C�"*��m���Ao��v �t4����eB���yIm��h�N%Ի���J=�{�����1��0+��?��ޏ��S�s�����׷Ln��OƎ���dN{0��-м�e�B �q�s��H��߼!)�QS�Kw}�皾e��we��0����Ev'�G膟� q�c*���A,���������%���( =m&�賮�a�<ݐ�)P�Ŧ�s^�d�XT�r�+�9�wB�;��>�~�v�km��à=B�*|�J�![�|&*7�To"�Yy	J�9DN�P�f)B,9@�w�}�c��t��+�����/H�e�Enk��y��2��X�	��>����7����6
�jU�F?	a��{]�?����^ޚ3�~�_�RZ!��g�� M�>�gt�|���{`���I�7����g���kl[:}�7��G%���\뗉Uk����*�j��N�mm��Vu��T�꯹���>>���B }p��z�@2,��x�KY���Y�h���% UUB�PL��������r�M��|�jev?mn\�����A�c
>�	�	���4k%���L����� �k1� �'��|��SMy�" �s��[��7��U�JY=�b�8�t�ŖWEz.�ʎ5;�a�8 ��������{�����v�ŵ]� C��?wx���S�K�-���oG7N�6'Ek��AJ�I�}��G�M�����j�y�l9 ���e���̱SRsX�6CC�'=fߤ���r�ߧϔ�jn?�Y�� �W��k����U��#	�s��ZJ�^Ǟ@�R���΍B!X	����6���L��޳�=�yxɊt�d�ZRMag�r_�*D�h���^E^��l���˲�s�_�A�Ϭ?��#����U�Q���ڽ&����^h�[M�8��:e�!�Bj�0��лV��y��{���,�i����lU�F�����s]� -�s%����4r%w9���^�������w�0�N�v�O�����T����wʨQ��	��}W^\`�2��4z�t=ż6�( ��e���W�/�POo]9��%���PrF�_�������Ҳ��ߦh}������/.cZzvE���6�a*�)X�E1y� uQ�������knـ�R�
��3���[��}d���5�fĥ(����k��@��'��mL4���u=����Æx��݉,��$�%��IƱF/�E����������b]9�F�:oY�}��Lh2�<L�&Q���$JyH��y�5���(�,��a��Z=��Q[��\}.�E��8���VK(0�Mո�kw^�yn�o~}�!R|тԋ��E�O��k��t|�JyR1p:���4�b���	_�0���<T�Gwِ$�'xὅ��:󭬒"��<�imʺ�dd��Q��Z��P����  ��6��n�Yb�5V��AO���*��F�B�w�n-t1�����̮����[Ϝ%G�k
$�o=+�?��Y���^��r�����kƖ�U�z��� PK   T��Zwxxz�  �  /   images/e78be1c6-81c8-4791-9ac1-5b77587554f8.png�wP�y��dm�����+*+�,/�DeiB�
".-�{`eW�PWC)
!���z�z�@@IHB����3wfg�{g�?����d�I~��;9�s���K��M��O ���kf� ` � ?9t��A����k�A p�}�)�����5��.�ϣ͊��d��l�ƳL�e���*R�>:=�e�(�!�<��|6��^���j���&��/�qC�D��=�ع9@�A����+Z�ⶵW��7��x߷Br���E�sh�@��},Κ���S�S�$*��;	q�qR�{�!��Ni,Q
;���'�qߙI&��D��B����8�>��I�p�, $��X6T5�^�`.�ɔ�wv�i6l�.qWNR���0�C ؖ�����p�2zכ�RBv%�G�Uٽy2�aI��3���:!�fw�	���2ݖď�#�%�z��#v_�Sl��%��#�H��l�b�W��7ӑR���}=ɱɆ�&'ZSG J��d�H���L{izq�[��Y��բ���[6յ��[m�$72i0sw���n;Q������ �J<QQ�Ts5[���0C��`b��@^��,��u���m��)��ٙ=ș^�S�0�.��ߦ9|ez�>����iZ��CG��Z����5!�0���RԴa+�r��������CV|�F%A��e���~������2c:��3t�����7G;��j8wC���;�@zz��d]�v=ˊ�����;�JF �l�Qֈ'JZ����}��2�h�!@B��݉=�{�:��֝��8���\�3=�P�C�
�vtPH�FB��K�L�fK4�\�|QCMȭ�_��w|>i����^����	|����ҬLT�I�"�tFK��xB�E��$�s3� �ż��q��n�
�
ďW|���#�AR$�+�Uu ���?)J�5�4�`��a�F��E>��t�����E�����3����[��V�Do5�H\kH�P�z=x�H��:o0���C�[��GϷn�t�Q���m+HP���K��G(�YaR��skB��f�?�X��~7Y2<6:���`�q�T��l�$SG>��\��&Dub<I庵���J��sp���g�"��vL��"��2�I��U���W8�!�FG�#���YgO�����oYq�!�K�<���H xkop6Rf����omp2� ʧ�� ��v�cs�S�ꚗ�%�b@ܝ���Z!��߉�b.�g��ϴv{!rZ[���Q 0�����iC�̝3E'��7��~�g͕Vo}��1N{<66�"3l���������r��n���l#���¬�&���;QF��[�?�>�aRP��E�Wp�1+����3���6�ن�����;����Z�ʈG�R]&��xF;
A(Ա���+}� ��-ש�!���zj���o�)7ى�o%Ö���i���U*tW���N�pDLiS�t��4<�_���u��w�ƫ�&=I5��h8٧�E�2S91ѪwS��r^���W�3<��6�O3�sg�f�6Z@:�������Ԑ��P^����)�f�����N>��N���� `#���\�+=��9YB�����;0G���ż��"�������/�^��d�����;�#���R\-Z��az�{u�q~��p ���\�u����L�eD���	W��D��bm�*����$�3Y��~���	�vGW���K��^K���:(�-޺0VFo��e��τN���z��S��x0��kc���"����J��!�jZ,����6|�5Ԩ�*W0ax��h������/�1��r�q'��ȫ-Ƭ�A�)�<q�G�84n�M	��h�#|��*��_�?�XB����@4�i9���	SK���:e������ٹ�%	�O�cc��NYǜ�U�����a�ۖ����-e7.$A�����֣�^��Uky����QJ���� H��L6��G�[���:�3***�~jаC7���@�~"F��uo�$��._�>XȄ!3��~+͘C�e��AV!��d��F��oPℏ&��+s�Ŏg� ����>��f��ȧ���#@�DQn���h �A���7ui�F�9��(I��=>6�����\���2�WO�;}Ǉ�]��8���c�볦��1'��i�ʧA��ażc�^�G�:�ڶK�Hſ��8�*�sm[\Rra��5�K)��Y���`�^���-uuZ����L��aF&QQ�R������G�ʤ�o�&h7���3YjH�յ���el�����i��śy�^1���[j 
``�v��2�.��2��'�ܙ�ٿ%��p8�����Q�(�AR�Uz����s�������7{�)Q��z焽����72p���*��k7K�M.�*�����k�G>m<&ꩵq��ppQ��m�̜���t�wVwoO��:V�e���Q�e�*P�^� �阹ؙ&�1������F���J�\Z��9��2F&��H/�����I��8!j�H�9�Жq���!�x}x�@[T�m�[���<�G�µ't��m���󸄡���q� �o��]�+]F��-��F|f$*�K�U)xVO�)����\�u�
��l��g8X�C\#�9t�'��p0���q�/{g^,�q�sO=���������rX��i�h�P����6s�%&E��I�CC;x,��ӋVI1�I/|*����d9#}&)V ���_�3B$��Nb�ճ���w��;��^y�����Ò���R�h��3�uu�K�e?������������������%�1������ָ��f�4l!�"�h��I� -`N��q�"-L���{sb�K!�T9�,x�Gd�}�,c愇zsͩ9<��(�-^���o|�-$���FƸ�"�M���E��
s)؉N�0�f�Rn���d�9B'$��O�dKզ����|�y����u:��Q�.��e��J덋�=��<;;��lu��j0;�)��f�lh,��;YۓSE?U-��x�j28�Mh�`���Ny�S Q��VEP.6ZX�l:����2!!!B���p���s�y�v�����
��w�?$L��*H�ƾL�0�����g^�Đ�D$�˛U&OC�ѕN5���.���'�v:�Z���� �q���tԀc1Eg!���T:�EmVb�~�� ���d2wձ���,�Խ� ��b+�N�����Ι���&
�~ɭK�|Fug�`w���:���""�*�ä�L";Ny�ǋ;%V;�#.�zXwi�h��ݏ�.�&����(���K��>]�?��$Y ��$��Z���x�"q�X�z�^�Rd����փ��x��ː�C5�,��7�蝯=���gv7_�A� 
0��L�.b���s�~~~�'�ڜ���W/�5��с�\�-���B�"�ͣa�SS����XFj�#�@��[p�a��!�(�n�p�����h���1J�M�L?� ҋ"n;W@.���'>[�W"�н���i��_�2��LַYe/P핯F�i4z,*#	vH���U��^k���:��޾�G@;��_�1i�Z��Ϻ�3_��ݾD��V�cQ�U���w�������
��Z��\�ׄ6u����E=�=�gXYƭ�7�`U�� I�>Tj�=��BaK�p�R�36:x{�N��5#-�;�<�/�:8X�6QE3Xo;@<huz��m��	��Z�T������2p�pxz7��,����A�1�=�.a���ӽ���9��ڱ/6���_�P�q�Ng�meD�1b^�nD����/6�P%�R.��%Rrk��@�6\Z�f��vжa�w yXYYYHU@�;�5|��g��rnC�S�.8�Fn���� ���OЯ��T�\N	[rX�!)�cB15��� �]{�Z�]d���B@�L���7��[Ix|@S���K��B�I��Vz䗀��� Dj�hӊ���)��*����A�+��+?σ�JL����J��:	�s��S�u)����[\a��.*))�5~0T(���",
��+|��B�k�0���וbgt�Ӡ��b�����S�i`H�|"F�����44��b2,���=���O�|��W���qs���x/��N-Mf<'���~�zm_�l��w��,�	�= ء��`������M��dEC�Q<8[�K��}�`7��w����v��ڬ�Oʖc?^T�p���H��II޻���Y�%$�H���Z���D�,���1��_����IHhPK��jqs��[\[)o�D���'P��<�-��;��,���؜�3��5^=p6&{#s���_���8^f��pJc�2��ܚ�=\�0����[w_$��$&�Ì�չ;�����э��<����Ι�ۘ�k����H�K]e�'=���:�]��js4,���	Ԓ�P����6ⷉK��[;��v��j�V��ػ�<�.�T�M�5	�X#���|+���l0jX��(=(P!32c��ؓ`��yxQ/<�y�J(��8D*�EEua�~)�!�|{�ɲ�S����R�|��o�8&�%��" 
�Ɥ�\6H!\�K*W<��l�I��Q3����Te���*�'k݊�	{�0.d'���ǅ�$,�a+�~�
�SK����cS��i��Zā©9e�C[^5��}@a�?����+���lGm��}Q'=�{ ��n~�s�G�PK   T��Z�+�s;  z;  /   images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngz;�ĉPNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ;IDATx��}�dU����z�B��=��ff��a� E��~���bXu]W�[]W�.:,b �H�!ϐ����=�=�su����ι�UuU�V�ou�Ztͭ���{���p�S^i���6���-��d~���q����n�%�c)E�Q��m2i�΅��Xi2S,��'m��.�FQ���-���Tm�����b0s�;B�~����e�>'Ax���;hW��������߾Om�P�-����sC�z�C�"�"�ZȐ4]PR
��m����5�������(|��D�>u�
e�ڶi2O]�m��$��0���9@m�������+��XҰд�OP�1,�|��� ��r�:�P�����:駙9E�)�3��5Pn�H��~{����mַ_��|���O[�)�٩����~qme����
`q���eIm�ō��!-o��/@Zє��7�dڶ}�|���m�
��-��!��he��x��u��6�o��~������_�$�.Z|��/LW����yf�!������o���h}/�|s�o5$��`qQ�)^�Z�,�̲��n�V4��8Ǧ=�`���e��J4#f4���`ZNѵ�iM4�h�Ry@��Y��3XL��Ч-F�����k6���,��LW���a:U��!�����
�<�.�0�x��N詔<�Q.�f�dw@���H�t5�C?z�v�f�ॕ�g(x����sYRa��]�^��Π�)�Ѡ�fF�Y�o0��C0��+p!�h�Iv;�H�8]���՗
 ڟ��h�4#��H���A<v����A2ɫe�{��caV(�(�Qiy����X����3�W3��@X��?�EI4c��j!]�"�� ,d}�D׮[涯�xSԥ
�3�2�b.CZrbe,�2i#;}Ƞ6�d5k��x�X�F�`��h�o\i:㼹�o�K/<��4�Mc6�*�Y1�g�b�)�L��E��>y�يܺ�652�=/�P�mWHa���H� M��Z
3�3B�����h'K*Mk1\��cC(?z of���.j�X�d�X/�Y�Ҽ���n��iE���1kD�͊��u'�_Q���n8��c�n0e��ym�à]2��ߊ�T�u��=��,�~O;�;=�K�n�"V�G�VB�zR��GV��D�q�[�Y��[.-n���Y� M���1�%B��Y�R3���������Ĳ&X)��X�X)\N���8��������{~���*��X��4#��j藃B�dY֓�P�6�t�H�����f�̥��>�Į�M<�U?!���|�}˜϶ؙ��<�����6��p҂���nz(CT��>���]���߲����[�D�چD".�a�.�߇v3"�8!iU��[ݼ��4j�9����#�x귏����c�觕o,}~�1��WRʂ܈�4�m���$/Ȑ1�6�������ӏ?��J1ޱ��,�u"1":���L��qO�Ik�Ѯ�!:�PuY1��+#1T66b� �x��)�E�z��P���ebJ�p!�BMQY5�=�@_��y����s1��҃ŭ��՚-�]��}��`�Lc�4�E1�8�hV҇6{F�+aAMezN��J�Lo�$�]]���u%P3,�)�c�D&����&�������D��ٝV�J���54���[`�B��2f�V;m-k5�uz0�?.�d��8M3ᯮ��ӅvR��OΨ�l^����C�3���'�(�Hf��,�o�&�^�n�^y�;_�n5m��F<���*�d�[�8��z`��J�`_��D��;��!��VRן,s���@g��p8PQQ!��O��eg�����)Y(��;��o�.X����ΚfX��0x	����k]#�k!;w#�3�:넥PK�C�`���:�E���=S\\�?���H*�Z���Ls�K&��H�h%h]ؾ�!<���(00�L*-�|1q50	}�82� ���X�N����o~�
�;C��W��";f�A�Ě�O���P�a�>2u�R*QP�c+t{0��|r(�F����f�ʈ�g6�^3܇�ۿV[�\d)n���e������Շ�o�C~4�r��U$���i�%I�T���좉�!��:aŮ#�#��Q�%e�����E���}Q�����<�h����4GؿEE"qv�ˎ3��B �%s�%�/- �3s��lᕖ`+�f=+��i�\f����P�I�ξ6}��-v~:����-�CH�&�|���{&Q�b%�z{�EgY�:����:������m�ɫ:��x�x�w�'���]�ǡ�*�t|�܍k�����F�UR`��K<��[0����o��zW�>QgGR�����'ahC�=�ъZ����Qd"���z��ƞy	�?7	�Q2��C&6������ߠ��sz�p����.���HX�2q~>����Iv�2ы�Ƣ/�'��g��iH�;}U�V�
��t�H��)�����0r3C�0������$��̶<p)�m�o�9hi�HN0>{Y�����E��CB�i|��jH6R}'�����4A�kj�*L���V^)�(��a���O��@�k٢�$��5@'"9������D°R{=Grt �8�d��Zh�{��TYEmbЏ����*�4�3�K�ӥzV�Ok_h�� �B�A�C�n��g�gƆ�coB��Y�����j�7�L�����	�W�L�c�]O���m�.[����u��P򳏣���a)��؝�G���!����|U�y��ct��H�1$b���gP���g2��?���J�$������-����v���'�p=���^��@/��%p�{���;܏�+އT�a��䋯��Ӆ���,�u�QMe]���G����:
^�!=Ǡ���#���,�C�����X�H�UP�e�p����lM`5w�.\.�f
7N:;(�*e�I��I#�JqzR�}�t��S��B�ij�V�DM�O�����]�@�O�~S�Q�-�
_K�*�O��Y/�Eu�?�pԏ�6�c1�%��t�sa<�l)�bvH�woC�?��.+��4�.�i�ҎE�J�5��@Z���"�=��Ϡ�̷kl4�IHU.���v��t�LP^�R� �i�T����5H�hB�:!���	!XH�����-��ό�BO&��0��#6��C���T����a�R����Ӣ��	Ȓ�>Mb��!{�P��nc�)�,>3$2��i�fxኘ�0(Ғ:Ns;q��C!��yU���S�c�7����k"@3 ��4�ii3S�y�Nz�J�X��e	v�"`�;���:�B��
A0-A��;��7"��FJ��H�B%]1y�� ��Ĩ(\OO�c�G���DL��J�[�x&�M0I�F�X�'��oC���n�`�D��L���H��hZ��	�}$@D�т�1��y����|4J$#~��I%��f�"ZS��� >�>��UM����f����v�_Nm��5<��`�D�'�UX���H��~*�#�l��*����C�o<uJ!fRC��0�K�����Y���ob�F����cV��?�=�x��&��e�~��%=
3#��U^�:���ue�8�)"��9�"��b\�~9��������i����7�?D�_nw��M�L/��M��s���s��9;d�P�=�O8V-2Z�du/FN ��_/�ȱ!�0՞v��}���%Bm��ϬϨ�0�zF�N��GF7��r�i[8](�X��uE�������$�����O~�n9c7]������Ӷ#��au�浈%�L�o�Z�E�$&�7�N�Y][��HN[��� 95�W_��	��c,>�N��w�����n�yYhln�燈����k���Mm��a�/&�Y�q=�B�lFt��z�G���0�g��9�^���f��� �iaC����!۬8���9h��=p8��$@�
��h��K������o����VU��uo�R��[i)DШ��d"���
�k4{�f����@����Ց4	�z��ڲ�O�'�E@����MŨM�\�v���k�ꢬ��xt0���T�(!�p�ظ}��CH�;�g�����,����K���Yh���!�ӱ��t� �L"M%�CX�*o>�?��C�y�dt6�����ק����g����eE�>-���/������x�p$f�8����ԑ� ���Ț�!�+��	��ʜv�=Dv����N�|�KA���7�B�1)�ljNQ}�=��;d�!�H���3��=���@s$�K�feD�f�C$FL/ll��;����V�<��7#�XN2�˕v2jB�˝�@�����D��k:��߷dt=Nl�p��\�5&�tQ%{|S��3C�sP� Ms�Éd<1�������d,mY��7�wS�_�wi�w�4��~�~0������Oi�Y4L���%�00HD�&R�F;�s�"����*��;�}���e����v���'F����f�&�_}��}�:�Ēp��������n�IcwN���:�r2����l=��X�픭��２�����׊>؅�������쇢1d����1r�LzA#���(�"�P�u�[�!,���сa������rܰe�	?��r�B;�Ey��a9�t�cU�;ػހ�؎��!A#�$��meY��s�5@����2$�	bH�]2�t�1c����\=�	v�����;��=32$�}n��a��ײ��}q�"��8��
�{��@������1V��@�4'8Dk���o���",;��-ȹz�����:�A~��ާ龳�!|����v�a�/ːI٭�myF�$��bV����b��w����A1CF3Sǿ����
s�'��?%|O�Oe*?v��fq��e3����-4���F{���>���^�f�_�������2�nN&S��=��b�,1�E�����F�B��b��n�Ӥ/��a���r�v�z&^Vp2\�2�'Ơ%�0Ek���ԊL$�����Y��U�����@g�^���#�u��{��뀕���2�#ƭ,J�}Ub�����R�B�׳�a��HRȯ��"���J���$�����
C_�sti��2-9$�)��UX��k��D��vH�D�}��C�"r
e�\���F�H�����.F���_q5��
��m@��qq��K�@���&�x2g��E��h�_��I�\04W)�Vݢ��(�{(�� �~qY��y�~�5(�{ 0=��`��P���pd4��ë��ِrb�x�LJ��W�vHn��gZ���Đ�e5,En��ȁ��\�$¿���h�I�7�#nm?�e�����]t����!�~z?�'3��hVL��(+�'�'�![&�Q�����PgL�f��~��AKP�@.f�Ёي6[��\�~Y��� ��K��ٞ"�'q�z����Bv:Qt�F���?���W��l%2�\3�r*��������)l�횋��&
�b�|6��٢������I�e2��8�W�2)5�XA.dk�������0���,>�\�[�b�W�@:�l�Ӫ�8�!C�.��]P|%P#!�D0�³(�~�����
{0�QKƌQҴI_�@xYhN4�0��� �(%�BɆ�z��"Y��j\ͫ���#��+p4��:�t��u#?���V��?�A��v��(m���b���#(��5��p��'VW��?$¶��8����Dp��g!�櫰U׊	ȓ�VY%Dw��A�ܙ0� ����m�VQE�"7��ar��L�@WS�@FB�Zb$$Y�s��1A�Ǎ�l�8w޿�E37N�1	 �z�D���C��XfxXYXD�XQ��fأ��Ӌ������G&M���`	b�ٽ��	�[��i'��:Խ�dB�GM��ޤ6g	z�{�i��썶��iO�<t@(��Ѐ�<�N#������V�
���;���$���[X:�z�ɈP��(�w͜La1�Ngo#�#@���pVz�a�Y��ٵ���2�cN�هk7��F��wb����U����H��B+�1�� �1%�oG���D�o�V��.�/��s�a�0_�
�e���3�Z����d��ayE3"yi�y�V��AݎǬn4�^��[����E�"�cq?~/��2:;;c�_V���w�Ia��~<m��Q|݇�#�X>�vZ��|�k_�/cC��=�1�G�B7�T,��A��r(ⓗ�gl�ǯ�n�:&,Di#��L�W�G�n���?�{�)���"Z �a�i��amA����Ah4I���'�4��p䅃�R�(�P,L�J�*�|�g�A<V�̄��-�i),�憢-`e��f������^�+.�^"\6��g������><�������L�1�q��V=����i��W�{��N�����&Y]L���$2v��D�B����C��'�Z�] ��
;Rezv�W��-H?|nR��6!nu�%{�T8��=�뗠{Z!�H@=F��ƿ��+�<�V5��	�3*I�S<�[u��ۧ݊+;����DҒ�2�� �ǘ�@~G1�~��P�?���9Kt8S1�w���x�[��~��⋌|�drF[�ۍ�r����b�)fw	�X�f�Kb,��C���aܶE��c/l�r��c>�b����!��C�¦�{�|��HZ�yb��V��p�57N#}L+��9,��}R'��>$��ܷ�����k�M������ʍh��M��'0�ė���-���3O}�8�u�pa8�"1�����%m�`.�p=3���'oڄ"~�9h�h�ӆ�n���>M�L�q�	����$��_R!]��5lw([�>4��<#'�K���6v�JvY�hʆ��
��꩘^6��>J����U��'�)�$%Oޓ"�y�Wx`�bC�V��eZ9�2��-�W^u��\�(Y@��сM��b�E��х�9�f��!M�C����ڇ����a�V�qZ���c�A8�[HIy��@�	B�_�S^J�,C3K�Y�E+��bS eǓm/f�*$�����6��d;_l�r] y!��?!�0����g�M��9�4pk;w ��DG�+~���tE#}�o��+j��	�� �(p�%^C�=.�Sߘ<�@�Y7Ŕߡh�W�ؐ���%
B_��͹�"[�Ղ��}E4�{C|���p�Q�dВ1X\ޜ��=�(j�:�&�XYY)`��~���	/��"�2CfIr���`E� ���F��w���;9����p(�7P7N��,%���ɺ��pVT�}�K-�U�\�>��Ŝ���0;6	�{��%dx}��_b�m/�ɑc�����,8�>I�e���R#1����*w�\(++CMu�	j��̙���ƻW�p�d�$�h�����'�R(�x�ڍ� a�A�rF����ņ���`�ß�{��<�JL�~�= _x"0�
N"�ԣ�#_DQ8���/��D�\9�+#!�]�E�2��.��d���
��p8��H���c�/ Or�I[,EQ���x�C�#�#�%��=�Xk��bt�0c������5t�n�v䈱`��K0U��g&̸'��tc�3��D��|����(��:Ay$�e��хzlJ+�EO���a�H�����pCQ,S[60�i@D�0Y�G��!f��8󯺺5U����#����h����Ç�q��֬�v1��*2��xb���21&���o3�~�, ���֞��}�8�2+�زb/J<L�4<<Hv��N��*n�?X��"�,p��!UUU���LQ$=I�B]�BkɴL�k�	��-R'(��D"�λ�����+�PRչ���l�%.�,���B3���hoG�"C�|[+�o-��V�sX���&e0���{:�%��԰̜?3z�V�ɑQ\�e+"�Q2��ˮ�h_m�ˠ0[U#G��{��̲"]ŵ��7^Ƿ�������[��pS�EL���FaUk�1����ۈ��|I@� [�Ծ��ń�M���[n)@YYg�0������,1��Ċ�8ғC`��۲
�S����E:�B�Dn'��GM3�FY4.�ˍ�d���Uը��Ĭ8���	�&�U���f��b�J7?���d�󷏡`7\֮]+c�I����}xf�s(&��,�l��l�㍞�4�5��e���@g�S"��}Y�#X��0���(��*����`���;	�T��d.I��4��@� ��P��]������8����F�57>�������>E�8�����Lx���!�Z�
M�a=�H�����µRc�#u�PS4�Uh�i-z������/��T���F��~�`��b�ϋ4d`` c��|�=Z׬1|\s0�Y�q�Dx�wX-� A���7�N�I���	T�!�h&O�m��+�*��[s)uj;��Иe�p�Y%%�������8�����~�H@�0S��q>��=�^{F��`k��\B bU�z�n����@U]����
l�Q�����"�W*.���D�*u����&h��D�z���3W��4F:�	x�⢘|ԟe�n����*�X%iى�{�xz8G�*HӺ��j�n���2�/L�"�Yb���8�&�M/̈��^�S�I[�I���ҁ�"SXI��e�S3F:�}�#���	|M9M�O{��]��4S�؞K�еե��|~���9��4�	�zpa�	����:��'�Q�NzM���l������.f�[IR�$�.�����!�zc^��Z�
Ȭ��ŃH��%f�[Ҁ6��Z"^��Ļ�}�S�np�EƲL7��PL6�H&�Ԝn�̭��s��%9����"�W"�����>�n�B�m�&l�&��<Y%�c��/��ƅ$}�<76���ǡ�3��7�� �Ua�I�����~�N6��[�R��a�<�^	��):�O��}8j+B�KAM���(F�:�*m9^�n'n�����p�ھ����Ӄ&E���2�W#zp�'���ߋ��h��ۍ`�	|��# ?��ag�x��Fr'!\'G�n>�p�x��L�-
��FFFP�~-���j�oWz!�IhW0~��aTUV���6��MU��?���M�Aó����7X�В��t�3���>�I��`�-��a��j���c�h.;����a�:Y��e�Wxx?�������=d�0�a8���|�)A�އ{t'A͙��YtG��Q�i"
;;N��|@A�P&��:E�IG�<St�2��|4>��b:A�k@(�0��DC��**��r/!}�z��ć�,Q����O�O���&K}�=��1?�)��p�s������y�#�8A+㹗;e�w;Ĕ���G04�4 Y͹]�*xq��Z��>.ғ\�Z=|P�K�rx9��l�_ºj%��<���ݹ�!|E�D���"��Jp�����&{g��{��9��� w[{��}��dk:�O�'��
�A���A�P19�uB��đ+pP��JJJP[[+���ȉ�jG�E6�<��|���R���&�1*�d����OJ�.H�z�
]$�͟��̨&��!�:Ja8hL~�����;}�L~?�L��3�!��8qa�'w�Y6��#�����_Ax�F��4�������L4�e�턪&V��k��N����Alڸ�_v�ܱ�>�(���66`���@��.�9b�X}%�^?��W�QRQm�(
�$<�.!㩟�ub�h*���j�e���+���#�����\e�����E"�|�>LsJ�M�c/��.,��`I���C�xP�_�au"�X<dHB3�Kl#�"�;���՝��34�Pz9M�Ёɭ�D��Kn�-[�o����.l�$�b����[�ك�^Z���G��P�����=�z��`��M��T�JZ����N$o5:6�[O���}b_���+Ѵ��h�x�U�2����=e;��,�d�`Ög���[C��~�$I݆h �FZ�	}3y�\YfH�~��L��$N�<�#�w=�����Σ����w�p�͂<�椩�oooǦ�N��%�}��b�5]�ޯ�iSv�p=�ů�g�^{�G��}�qU�r,�4�e�d6C��T��6�uB������'D���&�E6���14�M�P�#�1��*���g����fiqĐ�-�səL�����	#���iF�S6�['tF2�p9{���c�Qݼr�V���C���x&����g�_��ݮ���\�"T3��=b�o�8˫q4���چP,�DA�a�l4�W+	\alR��#d9��������:>t@���"�Y٧zc7���jY���Qw�����8����w
Ĕ�;Q���Rz�%����V��N�(Ny��{�J�uv��!v�gl�"�w2��+?���"�/kF�nZF��>�Bg��\�ؽ�m'��ϻ�x�`�F����� j�����
�9=ة{jjs��J7-�GFe@1^8A-i�1x_��&�1-��3�5�l=KlSQL>�4<��F�����M$F,(jY�T_����G2)n�8�H��@O���#�ۀ�@|g���+ϋ�
����!nK�Y&E޸|�����>�gt����Ҟ�獻�%��J��)���g���:Z��Hϓ�i#��X��o�.i�Wu<��,������蓄�톯_2��L���[$sv�M:jz*0�\�;׵""�<>��\,E�[o�,� C=��C����aD��`�!��@"��BǏ�H�y"P7���u?�G��pM ��S�˼�e���Fq�v.Ab�cɮ.���n#��!+���6\�!�^���$&�T1ƤQ�;t�C��=C4=��+���QxRQaq�R�s���=�:'iZ���[�l�d섽�A������u(�����dMK��J2�q�1b^�9����Ȟ�#�W����Қ�:q�
�q��%��O$MM�ά��i���x� ���	z�]n��WP�U���v$����b��P �w���%w<�˗§�IZ(�+T.ݶ��v}��O��b��^MR"J�]�+क�	؊��4{ݰON�E2:v�؎�&��(�B�f�N�׹�T�[OB���H���-kB�d��\�lTo1ĥ��2MԨ��1�Mے͓���0c�o~9p� .��,�P�n$��;O822��=>�.���J�:W�3!r`/�$�#���ZS�T$*�a:[�����!��4�Oı1��/�U�\���~��.x��Ι����v�vثV������?*�Qݼ =|5�����q�kP^���ŞF5F�՗s�#���{ϫ�QG��b�J�J��-^�3���J������*D{���E��R\����)	fV<����N������b�����"$߽[����w�}~�[σ�3���?������>�?R҄�n����)���	f����[�
S,���'1�%��r��r��mr�K<��r�6�S�y���c� 4;$�8X�<��� 0&i���?Ɨ��c��|���ouu��F�ܫp��X�Q���h"�,��+���z߻Cl�)�~´J�6��!!N����9
�(Ь����8c����/�燂�V��Õ��V�E�
����bqó�\A\�j���&�����w�,2��kk���l����ϣ%�%`�d��0�����!>�����y��D'�����w���s��>���p:��M����[��Zojj��3�YGɱ�����[k)�+�ov����Q>6������4����غ��<��X���-JHS'�H����Ŝ5<uޡ.�ϲ`�D;���`ǵ�@��Ni������POn�c~"C�H�ߣ-�{xX�>��?���ċ�}%#����
��8V�g�Y��8�ÿƱ�n|���ओNY�<Ax�d0�ǟ~/��Cv�W�ܣ͒�Ęs��/}5�ӳ;�����5��[��}��nNv��F'o��ྀ̽s�y���H�Q�;=����[}����H)(���o5�!��J��H�1�ɨ�Bh���0"�Bm_%��co�����W�2
�3�g����뱬��'wubt2A"vj�q���"S�"�p������GCC�4�]�������H�h�T%��&5Ǵ�[�DL�N�\V��V��kO�ˌC�/��T��N�J.��.��|1���nCI篰�p�8�)CW���KkE�n!���`�-��Ѩ084�~���wC�"]B�L���g�j��z�2�#�ܗ)ű�w@"�u*�0���7� ����2�f��ĔS��X�j� ��{L��s-湓�D4��]9�jxz�{F0H�т$=��컛&�
p{��Đ�׈�-�rbf�<x�o�ג�'S�֪
�%xxx�ؕ~୅�>H@`�.>���"�S���Hv���a��˅b�/3؉u��u�p�}⁹�����ԥ��V��Hb�}�rk������$#AB���1O5�����n!)Kbq��xN^�Yc0_�����Z*�X���l�t��!��.���^ ����rb�˛��ݐV4s���,^���&^��o=.H�{HR�y�Z��� ���9�u�J7�у��Z�hʐ��م�"ZeV���4�d`n�Ԍ5��3b�F��S��S�� ��E*?G���P������˦��=4�Q�ԧ�:D�w������01/.[�=0:�	������II�e����i!>�ה���5��$�1E3�2��դ�V\',vf}=��+�C]���!5��!J��o����^%^��o�.|}7�)%�'�@�h:�}�=��P�~9;��_A��ԋ[x�X"�X�J�����I!9����O[����@H��,����Ѹ�L$11a����,����pd҄G��IBN���"@F*G�,�XWg�{(,��܌6�y�t���Z-	�$�+��_�u]����Q��J�af�n�b�rb����Kj���̯�f��9V�"� ����@?�À֚��Nf$�)��03Z�u���{8���&ie�=D��_��H�S��Ey�6fF���A��/6�#qw�/g������z���p�l�ĺ�:���rPkYC�@asÝ�Ƥd�hξ`�7CK���O����<j�A2��Vd72�x�&o���k˪�%h�U�S���4.�[`#��&�z��T���*¦�H�z��[@c�j<.�pXr�}�b,	��������mB)zV��.�D��{Ǆ(.�C%=8��Wn9y-�����`Z�����eZ���gosh��R�MZ��!ۀ7�Z��;�$⪞J䗳kO�f����]QPJ��C𰴴T���WI��'�$���Cq+�	11øp�>��9�<���J�-ƓP]�VA�ׂ��W�U�}N�Q'�l�h�NXeS.��"��yC�@Y�?ہq\��f?�z������ET1�.o;k1Ђ�>CY5Ը�W�;V�-�O�<F�W�31�ҿh�2����}�����w��V��Ob��^�$��I7�����Dk��ܲn��د�DVn��n���K8W�&���w�Wހ�<⽯55�Ѽn\�R�߭��O+���B(k��k���r�D�-����)B5Y���G�[i���z�O߄3�p1ڡ����E�YMm%�VTQ8b����X�B*�� ;����I����,�Be^�'z�i����l����al�#��<�.흃�b����q����
�r(�t2t�3���Ca%[G�ض}ݍ��
.!yG�u=#�]����~X)��l��.o�U׊�B�3��S�.e�H�Npr��A��$�O�/Oo�K���P���	G���=�����xd2��[��U)A����C�2��e\���À3������$z��X�:q��d�P^b��t� ��G�f���V"�d��#�ә�+ԔP�)o����K���7�k�"�A��~�zACS���$ho�3�q���.~��KjX~/M��km�E�pޣwuؤ��c�W�V\0u��� ��IؿV>��V��SCp�+��2ـ�᰺G���BmGt�V���ŧ�,��&nk/rQۍh?8�J��S8�����ʋ�9m�� ���D�~"�l��E�E,�~R�c�e�H�ץ�Շ,�ʺ<4B�.#��M��&ɻI�3����Z���v�b�b�c$	4e�eR���5��}�m���~6Ĕ���^�i_���O��Ж��fb�&7y����c�g��$z�Ľ�ޏz��`����#�ȐcCLl�5N���ࣻ����bbV1��Lz��ڲ@R��3�1s[��m9�C�k+e?Sǜۈp�OL"�A"vS��2u�ܘ�D:� ���|.$��䤱?�&�B�L��mMNX/6��2F��ߊ����@5ι/���Ǡ�qz�S`9S�C D;FS���z��&fӜi?��|�-��?�
��m.BUg�h��AB�˃=�q�]x�tG��T�����q�\�I���e��c�i�xz�lgP��|���ݫ������� ��D��s�F��>z�7��Czl����`�&N8�','g�6�"�2��wb��;�hX.z��2V�|H��������>�H�A�h��]$����cF!CL�0��G��,Ѝ��^`�Wel�w?�'N�	[f�s�0C�$�rK�� D@�|Z�i7�9��8�ϫH)�%��a����A"f���B�4r��"��Ldm�=��OT�zf�qĬ,c���}�"�ħ��~3�x�
A�,����Z�U9���.��b?��SH�E<�h���"\��8�%���.�i$#p�*�"��
�E�!�sz�ԣ��	�=���d1QO�W��#�uςl�S�=��Y<�.D2���ȰnO{a�t͖���o�-\b�    IEND�B`�PK   T��Z��8�     /   images/fae81aff-08b8-4df9-bcc4-e5b22ddbe47f.png ���PNG

   IHDR   d   0   ��ߵ   	pHYs  �  ��+  �IDATx��{LGǿ����%��x>����#$4�V$��$bj�Hk�Gk��ӴFcSmRm��G��1M&���DC�P�b5ƴ����"��v�3�x�3���I~w{�������f�f%�Mww��#fo�v3+`v3+++�k�h]���1tA4�.����ゴ��`l�d�˾� tfU����@}�Q��f�OG���w�~Qz�}�e�xB"kd]�c�X	���4�l�`��p��)��&������A+�Β�7?�[D�����oS��'D8ȶ�s&�w?pݰ�M'�� ��q��%�z��Ճe6��2/��Y�b��݊P�!1��P!q���Dחfi�B�Aw��ܡ�(�Y؇���;Dc�6��DE��Ae�V^��6�|a�Nff���.&�/�13B��L��c�|:z�###>��="�b�9�i�$R���n�#�\��a�U�Xw�{\:��_Ҋ�p�\�^��W.ߜA)�(�S�|ǵ;��k���� %$3K�>k2z�L�=$%%q�40��H'��M�(����(	�[�M��/Lx8������*�R��؉1	�kt�>�DȒ��ڐ�	��B�d�@�[S���xꕏ_n�m��I�����ߧ^��RJc��!��Z�ZB�Wv�Y��p���h��G����$I�X�,�8RmQ���;��<�e�3�k���ʴ�������ӑ��	������Zf6^���ڵlTƏ���B^^JJJ���� h.�y9�E���|JKKa�Z�p[:�������M�6���MMM����C�׉J�\.�������u1�L���GZZ�����9��|����u.Jcc�*��#f9�f扉1?�(**���U
M�3\�=�8��p`bT���@mm�:���@YY�:��L��oh$�u��y*�%2�C�Q�u�.��?x������9؎g��᭖�ME��a!� ����d$·��w�ϟ���xP���c�!\�3x���J"w74�{������~�>䍆��n&F������Յ��Bu�X\\��P�z���#�����T477�#-Cx,џg�NL3���\tvv"''g�!�N�pA�0[���l^8'q���ߏӧO�#���VTVV�=$pAv����Xï�yK�yIHH����ՅN�S#N�.�W�Z�F	K�Rq�gpړ���l��4]��0Cz|���[+v�p����cBx����?�y���G� 
������N}�Z���٘����~�5���غ�!,�)L�Й����>	ǹ3Ȱ��
�O���������������kL�b���z�6�LU�J�`��Խ�,���_�/�=syY)_x���k�Ga�O�&\���(P��@�+ $9@L�R�{"���l��M���On�l/%U�R� .X�l�ޕ�v@ �#��}�B���������hB�lMaeL��ݦ.�N��N��x��l�h�2���������,,|!`��7�S�#���-i���[OB��{�	����������eK���x@}��D��	��i^GX�e˖�aܝ�nb�0�zncq_��Wʱ�
InOv}�TA��ڏ��GGu T �vv�����ס����PZ�1%�EJ����1>��<��GK�u&��1tA4�.����� �_�Vl�"pV>    IEND�B`�PK   T��Z��QZj  U?     jsons/user_defined.json�[�r�8���e�F�q��M��]�ė��Tm�R Ĭ�E���ɦ����E��8OK?ɔp����l�߆�יsW|L�Ϧ.����g�4|��pe�0�O����|��s�﫱ﰒ���}^�� -�0<��t���k2�X��E9�-���D�^O�n4��ǡH��\���@r��}Z}�NB�W�9vs[d�r5��뗙�ki�0(���C@!����s���S��|��	$�<�P�(��{�d�˹2�A�lz:�����p��?�泉�z�O�y��'
+�����ʿ��.@����f�a�����,���^� �g��βI5R%�#�F���B���d�����E<<,�E0�DW����{4�>����)�	�ӗ��[�7��>a4�TP9B"� S��FxR�g%�a�����������	d�Ю�y�n{.xBTlDI���>id�m\EK��~�� �7 �ʳUp Q�A��݀��1����6�_q�&�u'�h$R5"Ex�$�l�1�n��G�K`��Et;DM�$HF�4+ե�ZAAzKB��`�f���\������-v���5�`h1R]���`h� ڡr���JD04K�P��7u��o��o�������!1��|�2[��u�0_�Զ����iU.�ɢ����BXyH�r���w����Q~?۲W%�M6���m���bI��cժ��t�-Ų��R���M^�u0�C򩛖7�:;��O�]��U�1	'��wny��Eg�ZH��"�L�Ui8��|���E��!�l�)�n�5sT2c��!@1V@bC��ʄ�`�+?���(�V�A���	i�Hd%Q�-���`�zY����H�b	J�^c-����8*�W��++�� c;+�P_� ���*�\		��B$��@5�</�������7��*M:h�w���z�������u �	�����np������h�8�m��2���ă�
������Џ;�U�C�S�&{��&��u�� ]s4�S�C(8�WhC ��9h5�ܩ��h��{�v9O����^g(�����v���h���1͊G|ڄ���n��"�OHG����Gܑ���1�'�#�U���Ŗ�#�u���z'�x��.�.�<��<�b4��zP�v �
�5�����%�`�D�Z����餕Ja)I=����C\�Z����Ơ�����K���e� [vIv(�H��2�
�"��r>
Q>x�ؗH~�q��(�\R:��f��l��I�X�c��:����p�7znP�6esjpU!(��PS'	��kM���aG�QkkS\� ��;��L��5^�t������$T�e5�g���t�E��*z4ȦgS�?ˁ���=��If�����Y��g�����v~[�'W�L��[�B��GC?�fG[�;+�.��Xz2�Gj����|1M�F�����]�u[�.������"�*k�f�:sGA�|Z^g�uO& ��D��E���{M��i��	S1p>�4MS�ۉ�4'$�B/6�u��������s��^Ͻ�{=�z�����s��^Ͻ�{=���H�4����^�Yf�<L�,�����0���2
��
p"0`*�A�R%;�9fS( �Rj`
��W
;��� ����j���8����!��h���"x�e0������;j�������-<k��=�W���-�->�ur}�>���tÏ; �E���|�����G�c��n�aG�S�+p��E��`ˎ�<�l�[t�1�z7�M:}	.c�n���T��݀w��qX|�!�zG�#tpvq�|6|�)�EW�"|pvz�|*|�1^�7�<ypzs����@����ю�����e	T�.����f�����x�x����x<n����`������#c�9Q�xydT��Ԣێ�7���[T�Q���ȉ[4�Q�㫓���-��(Xr�rc[�9,���ߚ���j�VVɨ�����l�����f⺞�y7��(w�J�֕=�x��'�K�f�(�z`��^��(�z���˭�N��{�f\M��n��x�f���
��{6D�0d,�� ��,���i�^��U�����PK   T��Z����6  �R            ��    cirkitFile.jsonPK   T��Z����7  �  /           ���6  images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK   T��Zo�>��q  �q  /           ��3H  images/2cd737db-51bc-41eb-8762-f3273c40eae5.pngPK   T��ZFǫ�>  >  /           ��J�  images/3db32f6d-ca85-42a8-bb1f-49cf601f6ec4.pngPK   T��Z�Bʟ�� Y� /           ����  images/8b28e7b8-a93b-45a9-8e01-1e8c89928838.pngPK   T��ZN�v4	� m� /           ��� images/91e5cd07-2a88-4b0d-9128-72e2f992e16c.pngPK   T��Z�'k�  �  /           ���7 images/94f8244f-e118-4f93-ab30-835e0ca4f6e9.pngPK   T��Z�&�}[  y`  /           ��1O images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK   T��Z`$} [ /           ���� images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.pngPK   T��Z\���� �� /           ��a( images/c99f0c6d-affa-4fa1-a395-2aad1347a31a.pngPK   T��Zwxxz�  �  /           ���� images/e78be1c6-81c8-4791-9ac1-5b77587554f8.pngPK   T��Z�+�s;  z;  /           ���� images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngPK   T��Z��8�     /           ���% images/fae81aff-08b8-4df9-bcc4-e5b22ddbe47f.pngPK   T��Z��QZj  U?             ���, jsons/user_defined.jsonPK      �  �5   